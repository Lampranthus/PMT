library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity Test_LUT is
   port(
      CLK : in std_logic;
      I   : in  std_logic_vector(9 downto 0);
      A   : out std_logic_vector(17 downto 0)
      );
   end Test_LUT;

architecture ROM of Test_LUT is

subtype word_t is std_logic_vector(17 downto 0);
type memory_t is array(0 to 1023) of word_t;

signal rom : memory_t := (         -- Coefficient format 1.17
   "000000000000000000", -- Line 1   Column 1   Coefficient 0.00000000
   "010100100001111010", -- Line 1   Column 2   Coefficient 0.64155579
   "011010010110001010", -- Line 1   Column 3   Coefficient 0.82331848
   "010000010001011001", -- Line 1   Column 4   Coefficient 0.50849152
   "000010011111010011", -- Line 1   Column 5   Coefficient 0.07778168
   "111101011100010000", -- Line 1   Column 6   Coefficient -0.07995605
   "000001111101000010", -- Line 1   Column 7   Coefficient 0.06105042
   "000110101001101001", -- Line 1   Column 8   Coefficient 0.20783234
   "000011111011001101", -- Line 1   Column 9   Coefficient 0.12265778
   "111100100000110010", -- Line 1   Column 10   Coefficient -0.10899353
   "111001010001010000", -- Line 1   Column 11   Coefficient -0.21032715
   "111101100111011001", -- Line 1   Column 12   Coefficient -0.07451630
   "000010011111000101", -- Line 1   Column 13   Coefficient 0.07767487
   "111110001101000110", -- Line 1   Column 14   Coefficient -0.05610657
   "110000101101000011", -- Line 1   Column 15   Coefficient -0.47800446
   "100101111010100001", -- Line 1   Column 16   Coefficient -0.81517792
   "101010100001010101", -- Line 1   Column 17   Coefficient -0.67122650
   "111110011011100010", -- Line 1   Column 18   Coefficient -0.04905701
   "010011100000100111", -- Line 1   Column 19   Coefficient 0.60967255
   "011010100001111100", -- Line 1   Column 20   Coefficient 0.82907104
   "010001001110110001", -- Line 1   Column 21   Coefficient 0.53845978
   "000011001110011111", -- Line 1   Column 22   Coefficient 0.10082245
   "111101011010100101", -- Line 1   Column 23   Coefficient -0.08077240
   "000001100001011101", -- Line 1   Column 24   Coefficient 0.04758453
   "000110100010000111", -- Line 1   Column 25   Coefficient 0.20415497
   "000100010101101100", -- Line 1   Column 26   Coefficient 0.13558960
   "111100111110001000", -- Line 1   Column 27   Coefficient -0.09466553
   "111001001110100110", -- Line 1   Column 28   Coefficient -0.21162415
   "111101001100000010", -- Line 1   Column 29   Coefficient -0.08787537
   "000010010111100010", -- Line 1   Column 30   Coefficient 0.07398987
   "111110110110100001", -- Line 1   Column 31   Coefficient -0.03588104
   "110001101100001110", -- Line 1   Column 32   Coefficient -0.44715881
   "100110001111111001", -- Line 1   Column 33   Coefficient -0.80474091
   "101001101001010101", -- Line 1   Column 34   Coefficient -0.69857025
   "111100110111011011", -- Line 1   Column 35   Coefficient -0.09793854
   "010010011010111100", -- Line 1   Column 36   Coefficient 0.57565308
   "011010101000101100", -- Line 1   Column 37   Coefficient 0.83236694
   "010010001010110001", -- Line 1   Column 38   Coefficient 0.56775665
   "000100000000010101", -- Line 1   Column 39   Coefficient 0.12516022
   "111101011100000010", -- Line 1   Column 40   Coefficient -0.08006287
   "000001000110000110", -- Line 1   Column 41   Coefficient 0.03422546
   "000110011000010001", -- Line 1   Column 42   Coefficient 0.19934845
   "000100101110100001", -- Line 1   Column 43   Coefficient 0.14771271
   "111101011100101000", -- Line 1   Column 44   Coefficient -0.07977295
   "111001001110011100", -- Line 1   Column 45   Coefficient -0.21170044
   "111100110001001000", -- Line 1   Column 46   Coefficient -0.10101318
   "000010001101010010", -- Line 1   Column 47   Coefficient 0.06898499
   "111111011100110111", -- Line 1   Column 48   Coefficient -0.01715851
   "110010101011110101", -- Line 1   Column 49   Coefficient -0.41609955
   "100110101001110110", -- Line 1   Column 50   Coefficient -0.79206848
   "101000110110001101", -- Line 1   Column 51   Coefficient -0.72353363
   "111011010100000010", -- Line 1   Column 52   Coefficient -0.14646912
   "010001010001001001", -- Line 1   Column 53   Coefficient 0.53961945
   "011010101010010100", -- Line 1   Column 54   Coefficient 0.83316040
   "010011000101000110", -- Line 1   Column 55   Coefficient 0.59623718
   "000100110100101000", -- Line 1   Column 56   Coefficient 0.15069580
   "111101100000101100", -- Line 1   Column 57   Coefficient -0.07778931
   "000000101011001101", -- Line 1   Column 58   Coefficient 0.02109528
   "000110001100001010", -- Line 1   Column 59   Coefficient 0.19343567
   "000101000101100010", -- Line 1   Column 60   Coefficient 0.15895081
   "111101111100000110", -- Line 1   Column 61   Coefficient -0.06440735
   "111001010000110001", -- Line 1   Column 62   Coefficient -0.21056366
   "111100010110111001", -- Line 1   Column 63   Coefficient -0.11382294
   "000010000000011110", -- Line 1   Column 64   Coefficient 0.06272888
   "000000000000000000", -- Line 1   Column 65   Coefficient 0.00000000
   "110011101011100100", -- Line 1   Column 66   Coefficient -0.38497925
   "100111001000001001", -- Line 1   Column 67   Coefficient -0.77727509
   "101000001000001000", -- Line 1   Column 68   Coefficient -0.74603271
   "111001110001101111", -- Line 1   Column 69   Coefficient -0.19446564
   "010000000011011101", -- Line 1   Column 70   Coefficient 0.50168610
   "011010100110101101", -- Line 1   Column 71   Coefficient 0.83139801
   "010011111101011100", -- Line 1   Column 72   Coefficient 0.62374878
   "000101101011001011", -- Line 1   Column 73   Coefficient 0.17733002
   "111101101000101010", -- Line 1   Column 74   Coefficient -0.07389832
   "000000010000111111", -- Line 1   Column 75   Coefficient 0.00829315
   "000101111101111001", -- Line 1   Column 76   Coefficient 0.18647003
   "000101011010100111", -- Line 1   Column 77   Coefficient 0.16924286
   "111110011100011000", -- Line 1   Column 78   Coefficient -0.04864502
   "111001010101101000", -- Line 1   Column 79   Coefficient -0.20819092
   "111011111101100010", -- Line 1   Column 80   Coefficient -0.12620544
   "000001110001010001", -- Line 1   Column 81   Coefficient 0.05530548
   "000000011111110111", -- Line 1   Column 82   Coefficient 0.01555634
   "110100101011001000", -- Line 1   Column 83   Coefficient -0.35394287
   "100111101010100101", -- Line 1   Column 84   Coefficient -0.76045990
   "100111011111001101", -- Line 1   Column 85   Coefficient -0.76601410
   "111000010000111000", -- Line 1   Column 86   Coefficient -0.24176025
   "001110110010001000", -- Line 1   Column 87   Coefficient 0.46197510
   "011010011101110010", -- Line 1   Column 88   Coefficient 0.82704163
   "010100110011100000", -- Line 1   Column 89   Coefficient 0.65014648
   "000110100011110010", -- Line 1   Column 90   Coefficient 0.20497131
   "111101110011111111", -- Line 1   Column 91   Coefficient -0.06836700
   "111111110111101100", -- Line 1   Column 92   Coefficient -0.00405884
   "000101101101100110", -- Line 1   Column 93   Coefficient 0.17851257
   "000101101101100111", -- Line 1   Column 94   Coefficient 0.17852020
   "111110111101010000", -- Line 1   Column 95   Coefficient -0.03259277
   "111001011100111110", -- Line 1   Column 96   Coefficient -0.20460510
   "111011100101001111", -- Line 1   Column 97   Coefficient -0.13806915
   "000001011111110111", -- Line 1   Column 98   Coefficient 0.04680634
   "000000111100010110", -- Line 1   Column 99   Coefficient 0.02946472
   "110101101010001101", -- Line 1   Column 100   Coefficient -0.32314301
   "101000010000111100", -- Line 1   Column 101   Coefficient -0.74172974
   "100110111011100001", -- Line 1   Column 102   Coefficient -0.78343964
   "110110110001110010", -- Line 1   Column 103   Coefficient -0.28819275
   "001101011101011101", -- Line 1   Column 104   Coefficient 0.42063141
   "011010001111100001", -- Line 1   Column 105   Coefficient 0.82007599
   "010101100110111110", -- Line 1   Column 106   Coefficient 0.67527771
   "000111011110001100", -- Line 1   Column 107   Coefficient 0.23348999
   "111110000010101111", -- Line 1   Column 108   Coefficient -0.06116486
   "111111011111100010", -- Line 1   Column 109   Coefficient -0.01585388
   "000101011011011000", -- Line 1   Column 110   Coefficient 0.16961670
   "000101111110011101", -- Line 1   Column 111   Coefficient 0.18674469
   "111111011110100001", -- Line 1   Column 112   Coefficient -0.01634979
   "111001100110110001", -- Line 1   Column 113   Coefficient -0.19982147
   "111011001110001101", -- Line 1   Column 114   Coefficient -0.14931488
   "000001001100011101", -- Line 1   Column 115   Coefficient 0.03733063
   "000001010101011100", -- Line 1   Column 116   Coefficient 0.04171753
   "110110101000100010", -- Line 1   Column 117   Coefficient -0.29270935
   "101000111010111110", -- Line 1   Column 118   Coefficient -0.72120667
   "100110011101001001", -- Line 1   Column 119   Coefficient -0.79827118
   "110101010100110101", -- Line 1   Column 120   Coefficient -0.33358002
   "001100000101101101", -- Line 1   Column 121   Coefficient 0.37778473
   "011001111011111000", -- Line 1   Column 122   Coefficient 0.81048584
   "010110010111100101", -- Line 1   Column 123   Coefficient 0.69901276
   "001000011010001011", -- Line 1   Column 124   Coefficient 0.26277924
   "111110010100111011", -- Line 1   Column 125   Coefficient -0.05228424
   "111111001000101111", -- Line 1   Column 126   Coefficient -0.02698517
   "000101000111011001", -- Line 1   Column 127   Coefficient 0.15985870
   "000110001101000001", -- Line 1   Column 128   Coefficient 0.19385529
   "000000000000000000", -- Line 1   Column 129   Coefficient 0.00000000
   "111001110010111111", -- Line 1   Column 130   Coefficient -0.19385529
   "111010111000100111", -- Line 1   Column 131   Coefficient -0.15985870
   "000000110111010001", -- Line 1   Column 132   Coefficient 0.02698517
   "000001101011000101", -- Line 1   Column 133   Coefficient 0.05228424
   "110111100101110101", -- Line 1   Column 134   Coefficient -0.26277924
   "101001101000011011", -- Line 1   Column 135   Coefficient -0.69901276
   "100110000100001000", -- Line 1   Column 136   Coefficient -0.81048584
   "110011111010010011", -- Line 1   Column 137   Coefficient -0.37778473
   "001010101011001011", -- Line 1   Column 138   Coefficient 0.33358002
   "011001100010110111", -- Line 1   Column 139   Coefficient 0.79827118
   "010111000101000010", -- Line 1   Column 140   Coefficient 0.72120667
   "001001010111011110", -- Line 1   Column 141   Coefficient 0.29270935
   "111110101010100100", -- Line 1   Column 142   Coefficient -0.04171753
   "111110110011100011", -- Line 1   Column 143   Coefficient -0.03733063
   "000100110001110011", -- Line 1   Column 144   Coefficient 0.14931488
   "000110011001001111", -- Line 1   Column 145   Coefficient 0.19982147
   "000000100001011111", -- Line 1   Column 146   Coefficient 0.01634979
   "111010000001100011", -- Line 1   Column 147   Coefficient -0.18674469
   "111010100100101000", -- Line 1   Column 148   Coefficient -0.16961670
   "000000100000011110", -- Line 1   Column 149   Coefficient 0.01585388
   "000001111101010001", -- Line 1   Column 150   Coefficient 0.06116486
   "111000100001110100", -- Line 1   Column 151   Coefficient -0.23348999
   "101010011001000010", -- Line 1   Column 152   Coefficient -0.67527771
   "100101110000011111", -- Line 1   Column 153   Coefficient -0.82007599
   "110010100010100011", -- Line 1   Column 154   Coefficient -0.42063141
   "001001001110001110", -- Line 1   Column 155   Coefficient 0.28819275
   "011001000100011111", -- Line 1   Column 156   Coefficient 0.78343964
   "010111101111000100", -- Line 1   Column 157   Coefficient 0.74172974
   "001010010101110011", -- Line 1   Column 158   Coefficient 0.32314301
   "111111000011101010", -- Line 1   Column 159   Coefficient -0.02946472
   "111110100000001001", -- Line 1   Column 160   Coefficient -0.04680634
   "000100011010110001", -- Line 1   Column 161   Coefficient 0.13806915
   "000110100011000010", -- Line 1   Column 162   Coefficient 0.20460510
   "000001000010110000", -- Line 1   Column 163   Coefficient 0.03259277
   "111010010010011001", -- Line 1   Column 164   Coefficient -0.17852020
   "111010010010011010", -- Line 1   Column 165   Coefficient -0.17851257
   "000000001000010100", -- Line 1   Column 166   Coefficient 0.00405884
   "000010001100000001", -- Line 1   Column 167   Coefficient 0.06836700
   "111001011100001110", -- Line 1   Column 168   Coefficient -0.20497131
   "101011001100100000", -- Line 1   Column 169   Coefficient -0.65014648
   "100101100010001110", -- Line 1   Column 170   Coefficient -0.82704163
   "110001001101111000", -- Line 1   Column 171   Coefficient -0.46197510
   "000111101111001000", -- Line 1   Column 172   Coefficient 0.24176025
   "011000100000110011", -- Line 1   Column 173   Coefficient 0.76601410
   "011000010101011011", -- Line 1   Column 174   Coefficient 0.76045990
   "001011010100111000", -- Line 1   Column 175   Coefficient 0.35394287
   "111111100000001001", -- Line 1   Column 176   Coefficient -0.01555634
   "111110001110101111", -- Line 1   Column 177   Coefficient -0.05530548
   "000100000010011110", -- Line 1   Column 178   Coefficient 0.12620544
   "000110101010011000", -- Line 1   Column 179   Coefficient 0.20819092
   "000001100011101000", -- Line 1   Column 180   Coefficient 0.04864502
   "111010100101011001", -- Line 1   Column 181   Coefficient -0.16924286
   "111010000010000111", -- Line 1   Column 182   Coefficient -0.18647003
   "111111101111000001", -- Line 1   Column 183   Coefficient -0.00829315
   "000010010111010110", -- Line 1   Column 184   Coefficient 0.07389832
   "111010010100110101", -- Line 1   Column 185   Coefficient -0.17733002
   "101100000010100100", -- Line 1   Column 186   Coefficient -0.62374878
   "100101011001010011", -- Line 1   Column 187   Coefficient -0.83139801
   "101111111100100011", -- Line 1   Column 188   Coefficient -0.50168610
   "000110001110010001", -- Line 1   Column 189   Coefficient 0.19446564
   "010111110111111000", -- Line 1   Column 190   Coefficient 0.74603271
   "011000110111110111", -- Line 1   Column 191   Coefficient 0.77727509
   "001100010100011100", -- Line 1   Column 192   Coefficient 0.38497925
   "000000000000000000", -- Line 1   Column 193   Coefficient 0.00000000
   "111101111111100010", -- Line 1   Column 194   Coefficient -0.06272888
   "000011101001000111", -- Line 1   Column 195   Coefficient 0.11382294
   "000110101111001111", -- Line 1   Column 196   Coefficient 0.21056366
   "000010000011111010", -- Line 1   Column 197   Coefficient 0.06440735
   "111010111010011110", -- Line 1   Column 198   Coefficient -0.15895081
   "111001110011110110", -- Line 1   Column 199   Coefficient -0.19343567
   "111111010100110011", -- Line 1   Column 200   Coefficient -0.02109528
   "000010011111010100", -- Line 1   Column 201   Coefficient 0.07778931
   "111011001011011000", -- Line 1   Column 202   Coefficient -0.15069580
   "101100111010111010", -- Line 1   Column 203   Coefficient -0.59623718
   "100101010101101100", -- Line 1   Column 204   Coefficient -0.83316040
   "101110101110110111", -- Line 1   Column 205   Coefficient -0.53961945
   "000100101011111110", -- Line 1   Column 206   Coefficient 0.14646912
   "010111001001110011", -- Line 1   Column 207   Coefficient 0.72353363
   "011001010110001010", -- Line 1   Column 208   Coefficient 0.79206848
   "001101010100001011", -- Line 1   Column 209   Coefficient 0.41609955
   "000000100011001001", -- Line 1   Column 210   Coefficient 0.01715851
   "111101110010101110", -- Line 1   Column 211   Coefficient -0.06898499
   "000011001110111000", -- Line 1   Column 212   Coefficient 0.10101318
   "000110110001100100", -- Line 1   Column 213   Coefficient 0.21170044
   "000010100011011000", -- Line 1   Column 214   Coefficient 0.07977295
   "111011010001011111", -- Line 1   Column 215   Coefficient -0.14771271
   "111001100111101111", -- Line 1   Column 216   Coefficient -0.19934845
   "111110111001111010", -- Line 1   Column 217   Coefficient -0.03422546
   "000010100011111110", -- Line 1   Column 218   Coefficient 0.08006287
   "111011111111101011", -- Line 1   Column 219   Coefficient -0.12516022
   "101101110101001111", -- Line 1   Column 220   Coefficient -0.56775665
   "100101010111010100", -- Line 1   Column 221   Coefficient -0.83236694
   "101101100101000100", -- Line 1   Column 222   Coefficient -0.57565308
   "000011001000100101", -- Line 1   Column 223   Coefficient 0.09793854
   "010110010110101011", -- Line 1   Column 224   Coefficient 0.69857025
   "011001110000000111", -- Line 1   Column 225   Coefficient 0.80474091
   "001110010011110010", -- Line 1   Column 226   Coefficient 0.44715881
   "000001001001011111", -- Line 1   Column 227   Coefficient 0.03588104
   "111101101000011110", -- Line 1   Column 228   Coefficient -0.07398987
   "000010110011111110", -- Line 1   Column 229   Coefficient 0.08787537
   "000110110001011010", -- Line 1   Column 230   Coefficient 0.21162415
   "000011000001111000", -- Line 1   Column 231   Coefficient 0.09466553
   "111011101010010100", -- Line 1   Column 232   Coefficient -0.13558960
   "111001011101111001", -- Line 1   Column 233   Coefficient -0.20415497
   "111110011110100011", -- Line 1   Column 234   Coefficient -0.04758453
   "000010100101011011", -- Line 1   Column 235   Coefficient 0.08077240
   "111100110001100001", -- Line 1   Column 236   Coefficient -0.10082245
   "101110110001001111", -- Line 1   Column 237   Coefficient -0.53845978
   "100101011110000100", -- Line 1   Column 238   Coefficient -0.82907104
   "101100011111011001", -- Line 1   Column 239   Coefficient -0.60967255
   "000001100100011110", -- Line 1   Column 240   Coefficient 0.04905701
   "010101011110101011", -- Line 1   Column 241   Coefficient 0.67122650
   "011010000101011111", -- Line 1   Column 242   Coefficient 0.81517792
   "001111010010111101", -- Line 1   Column 243   Coefficient 0.47800446
   "000001110010111010", -- Line 1   Column 244   Coefficient 0.05610657
   "111101100000111011", -- Line 1   Column 245   Coefficient -0.07767487
   "000010011000100111", -- Line 1   Column 246   Coefficient 0.07451630
   "000110101110110000", -- Line 1   Column 247   Coefficient 0.21032715
   "000011011111001110", -- Line 1   Column 248   Coefficient 0.10899353
   "111100000100110011", -- Line 1   Column 249   Coefficient -0.12265778
   "111001010110010111", -- Line 1   Column 250   Coefficient -0.20783234
   "111110000010111110", -- Line 1   Column 251   Coefficient -0.06105042
   "000010100011110000", -- Line 1   Column 252   Coefficient 0.07995605
   "111101100000101101", -- Line 1   Column 253   Coefficient -0.07778168
   "101111101110100111", -- Line 1   Column 254   Coefficient -0.50849152
   "100101101001110110", -- Line 1   Column 255   Coefficient -0.82331848
   "101011011110000110", -- Line 1   Column 256   Coefficient -0.64155579
   "000000000000000000", -- Line 1   Column 257   Coefficient 0.00000000
   "010100100001111010", -- Line 1   Column 258   Coefficient 0.64155579
   "011010010110001010", -- Line 1   Column 259   Coefficient 0.82331848
   "010000010001011001", -- Line 1   Column 260   Coefficient 0.50849152
   "000010011111010011", -- Line 1   Column 261   Coefficient 0.07778168
   "111101011100010000", -- Line 1   Column 262   Coefficient -0.07995605
   "000001111101000010", -- Line 1   Column 263   Coefficient 0.06105042
   "000110101001101001", -- Line 1   Column 264   Coefficient 0.20783234
   "000011111011001101", -- Line 1   Column 265   Coefficient 0.12265778
   "111100100000110010", -- Line 1   Column 266   Coefficient -0.10899353
   "111001010001010000", -- Line 1   Column 267   Coefficient -0.21032715
   "111101100111011001", -- Line 1   Column 268   Coefficient -0.07451630
   "000010011111000101", -- Line 1   Column 269   Coefficient 0.07767487
   "111110001101000110", -- Line 1   Column 270   Coefficient -0.05610657
   "110000101101000011", -- Line 1   Column 271   Coefficient -0.47800446
   "100101111010100001", -- Line 1   Column 272   Coefficient -0.81517792
   "101010100001010101", -- Line 1   Column 273   Coefficient -0.67122650
   "111110011011100010", -- Line 1   Column 274   Coefficient -0.04905701
   "010011100000100111", -- Line 1   Column 275   Coefficient 0.60967255
   "011010100001111100", -- Line 1   Column 276   Coefficient 0.82907104
   "010001001110110001", -- Line 1   Column 277   Coefficient 0.53845978
   "000011001110011111", -- Line 1   Column 278   Coefficient 0.10082245
   "111101011010100101", -- Line 1   Column 279   Coefficient -0.08077240
   "000001100001011101", -- Line 1   Column 280   Coefficient 0.04758453
   "000110100010000111", -- Line 1   Column 281   Coefficient 0.20415497
   "000100010101101100", -- Line 1   Column 282   Coefficient 0.13558960
   "111100111110001000", -- Line 1   Column 283   Coefficient -0.09466553
   "111001001110100110", -- Line 1   Column 284   Coefficient -0.21162415
   "111101001100000010", -- Line 1   Column 285   Coefficient -0.08787537
   "000010010111100010", -- Line 1   Column 286   Coefficient 0.07398987
   "111110110110100001", -- Line 1   Column 287   Coefficient -0.03588104
   "110001101100001110", -- Line 1   Column 288   Coefficient -0.44715881
   "100110001111111001", -- Line 1   Column 289   Coefficient -0.80474091
   "101001101001010101", -- Line 1   Column 290   Coefficient -0.69857025
   "111100110111011011", -- Line 1   Column 291   Coefficient -0.09793854
   "010010011010111100", -- Line 1   Column 292   Coefficient 0.57565308
   "011010101000101100", -- Line 1   Column 293   Coefficient 0.83236694
   "010010001010110001", -- Line 1   Column 294   Coefficient 0.56775665
   "000100000000010101", -- Line 1   Column 295   Coefficient 0.12516022
   "111101011100000010", -- Line 1   Column 296   Coefficient -0.08006287
   "000001000110000110", -- Line 1   Column 297   Coefficient 0.03422546
   "000110011000010001", -- Line 1   Column 298   Coefficient 0.19934845
   "000100101110100001", -- Line 1   Column 299   Coefficient 0.14771271
   "111101011100101000", -- Line 1   Column 300   Coefficient -0.07977295
   "111001001110011100", -- Line 1   Column 301   Coefficient -0.21170044
   "111100110001001000", -- Line 1   Column 302   Coefficient -0.10101318
   "000010001101010010", -- Line 1   Column 303   Coefficient 0.06898499
   "111111011100110111", -- Line 1   Column 304   Coefficient -0.01715851
   "110010101011110101", -- Line 1   Column 305   Coefficient -0.41609955
   "100110101001110110", -- Line 1   Column 306   Coefficient -0.79206848
   "101000110110001101", -- Line 1   Column 307   Coefficient -0.72353363
   "111011010100000010", -- Line 1   Column 308   Coefficient -0.14646912
   "010001010001001001", -- Line 1   Column 309   Coefficient 0.53961945
   "011010101010010100", -- Line 1   Column 310   Coefficient 0.83316040
   "010011000101000110", -- Line 1   Column 311   Coefficient 0.59623718
   "000100110100101000", -- Line 1   Column 312   Coefficient 0.15069580
   "111101100000101100", -- Line 1   Column 313   Coefficient -0.07778931
   "000000101011001101", -- Line 1   Column 314   Coefficient 0.02109528
   "000110001100001010", -- Line 1   Column 315   Coefficient 0.19343567
   "000101000101100010", -- Line 1   Column 316   Coefficient 0.15895081
   "111101111100000110", -- Line 1   Column 317   Coefficient -0.06440735
   "111001010000110001", -- Line 1   Column 318   Coefficient -0.21056366
   "111100010110111001", -- Line 1   Column 319   Coefficient -0.11382294
   "000010000000011110", -- Line 1   Column 320   Coefficient 0.06272888
   "000000000000000000", -- Line 1   Column 321   Coefficient 0.00000000
   "110011101011100100", -- Line 1   Column 322   Coefficient -0.38497925
   "100111001000001001", -- Line 1   Column 323   Coefficient -0.77727509
   "101000001000001000", -- Line 1   Column 324   Coefficient -0.74603271
   "111001110001101111", -- Line 1   Column 325   Coefficient -0.19446564
   "010000000011011101", -- Line 1   Column 326   Coefficient 0.50168610
   "011010100110101101", -- Line 1   Column 327   Coefficient 0.83139801
   "010011111101011100", -- Line 1   Column 328   Coefficient 0.62374878
   "000101101011001011", -- Line 1   Column 329   Coefficient 0.17733002
   "111101101000101010", -- Line 1   Column 330   Coefficient -0.07389832
   "000000010000111111", -- Line 1   Column 331   Coefficient 0.00829315
   "000101111101111001", -- Line 1   Column 332   Coefficient 0.18647003
   "000101011010100111", -- Line 1   Column 333   Coefficient 0.16924286
   "111110011100011000", -- Line 1   Column 334   Coefficient -0.04864502
   "111001010101101000", -- Line 1   Column 335   Coefficient -0.20819092
   "111011111101100010", -- Line 1   Column 336   Coefficient -0.12620544
   "000001110001010001", -- Line 1   Column 337   Coefficient 0.05530548
   "000000011111110111", -- Line 1   Column 338   Coefficient 0.01555634
   "110100101011001000", -- Line 1   Column 339   Coefficient -0.35394287
   "100111101010100101", -- Line 1   Column 340   Coefficient -0.76045990
   "100111011111001101", -- Line 1   Column 341   Coefficient -0.76601410
   "111000010000111000", -- Line 1   Column 342   Coefficient -0.24176025
   "001110110010001000", -- Line 1   Column 343   Coefficient 0.46197510
   "011010011101110010", -- Line 1   Column 344   Coefficient 0.82704163
   "010100110011100000", -- Line 1   Column 345   Coefficient 0.65014648
   "000110100011110010", -- Line 1   Column 346   Coefficient 0.20497131
   "111101110011111111", -- Line 1   Column 347   Coefficient -0.06836700
   "111111110111101100", -- Line 1   Column 348   Coefficient -0.00405884
   "000101101101100110", -- Line 1   Column 349   Coefficient 0.17851257
   "000101101101100111", -- Line 1   Column 350   Coefficient 0.17852020
   "111110111101010000", -- Line 1   Column 351   Coefficient -0.03259277
   "111001011100111110", -- Line 1   Column 352   Coefficient -0.20460510
   "111011100101001111", -- Line 1   Column 353   Coefficient -0.13806915
   "000001011111110111", -- Line 1   Column 354   Coefficient 0.04680634
   "000000111100010110", -- Line 1   Column 355   Coefficient 0.02946472
   "110101101010001101", -- Line 1   Column 356   Coefficient -0.32314301
   "101000010000111100", -- Line 1   Column 357   Coefficient -0.74172974
   "100110111011100001", -- Line 1   Column 358   Coefficient -0.78343964
   "110110110001110010", -- Line 1   Column 359   Coefficient -0.28819275
   "001101011101011101", -- Line 1   Column 360   Coefficient 0.42063141
   "011010001111100001", -- Line 1   Column 361   Coefficient 0.82007599
   "010101100110111110", -- Line 1   Column 362   Coefficient 0.67527771
   "000111011110001100", -- Line 1   Column 363   Coefficient 0.23348999
   "111110000010101111", -- Line 1   Column 364   Coefficient -0.06116486
   "111111011111100010", -- Line 1   Column 365   Coefficient -0.01585388
   "000101011011011000", -- Line 1   Column 366   Coefficient 0.16961670
   "000101111110011101", -- Line 1   Column 367   Coefficient 0.18674469
   "111111011110100001", -- Line 1   Column 368   Coefficient -0.01634979
   "111001100110110001", -- Line 1   Column 369   Coefficient -0.19982147
   "111011001110001101", -- Line 1   Column 370   Coefficient -0.14931488
   "000001001100011101", -- Line 1   Column 371   Coefficient 0.03733063
   "000001010101011100", -- Line 1   Column 372   Coefficient 0.04171753
   "110110101000100010", -- Line 1   Column 373   Coefficient -0.29270935
   "101000111010111110", -- Line 1   Column 374   Coefficient -0.72120667
   "100110011101001001", -- Line 1   Column 375   Coefficient -0.79827118
   "110101010100110101", -- Line 1   Column 376   Coefficient -0.33358002
   "001100000101101101", -- Line 1   Column 377   Coefficient 0.37778473
   "011001111011111000", -- Line 1   Column 378   Coefficient 0.81048584
   "010110010111100101", -- Line 1   Column 379   Coefficient 0.69901276
   "001000011010001011", -- Line 1   Column 380   Coefficient 0.26277924
   "111110010100111011", -- Line 1   Column 381   Coefficient -0.05228424
   "111111001000101111", -- Line 1   Column 382   Coefficient -0.02698517
   "000101000111011001", -- Line 1   Column 383   Coefficient 0.15985870
   "000110001101000001", -- Line 1   Column 384   Coefficient 0.19385529
   "000000000000000000", -- Line 1   Column 385   Coefficient 0.00000000
   "111001110010111111", -- Line 1   Column 386   Coefficient -0.19385529
   "111010111000100111", -- Line 1   Column 387   Coefficient -0.15985870
   "000000110111010001", -- Line 1   Column 388   Coefficient 0.02698517
   "000001101011000101", -- Line 1   Column 389   Coefficient 0.05228424
   "110111100101110101", -- Line 1   Column 390   Coefficient -0.26277924
   "101001101000011011", -- Line 1   Column 391   Coefficient -0.69901276
   "100110000100001000", -- Line 1   Column 392   Coefficient -0.81048584
   "110011111010010011", -- Line 1   Column 393   Coefficient -0.37778473
   "001010101011001011", -- Line 1   Column 394   Coefficient 0.33358002
   "011001100010110111", -- Line 1   Column 395   Coefficient 0.79827118
   "010111000101000010", -- Line 1   Column 396   Coefficient 0.72120667
   "001001010111011110", -- Line 1   Column 397   Coefficient 0.29270935
   "111110101010100100", -- Line 1   Column 398   Coefficient -0.04171753
   "111110110011100011", -- Line 1   Column 399   Coefficient -0.03733063
   "000100110001110011", -- Line 1   Column 400   Coefficient 0.14931488
   "000110011001001111", -- Line 1   Column 401   Coefficient 0.19982147
   "000000100001011111", -- Line 1   Column 402   Coefficient 0.01634979
   "111010000001100011", -- Line 1   Column 403   Coefficient -0.18674469
   "111010100100101000", -- Line 1   Column 404   Coefficient -0.16961670
   "000000100000011110", -- Line 1   Column 405   Coefficient 0.01585388
   "000001111101010001", -- Line 1   Column 406   Coefficient 0.06116486
   "111000100001110100", -- Line 1   Column 407   Coefficient -0.23348999
   "101010011001000010", -- Line 1   Column 408   Coefficient -0.67527771
   "100101110000011111", -- Line 1   Column 409   Coefficient -0.82007599
   "110010100010100011", -- Line 1   Column 410   Coefficient -0.42063141
   "001001001110001110", -- Line 1   Column 411   Coefficient 0.28819275
   "011001000100011111", -- Line 1   Column 412   Coefficient 0.78343964
   "010111101111000100", -- Line 1   Column 413   Coefficient 0.74172974
   "001010010101110011", -- Line 1   Column 414   Coefficient 0.32314301
   "111111000011101010", -- Line 1   Column 415   Coefficient -0.02946472
   "111110100000001001", -- Line 1   Column 416   Coefficient -0.04680634
   "000100011010110001", -- Line 1   Column 417   Coefficient 0.13806915
   "000110100011000010", -- Line 1   Column 418   Coefficient 0.20460510
   "000001000010110000", -- Line 1   Column 419   Coefficient 0.03259277
   "111010010010011001", -- Line 1   Column 420   Coefficient -0.17852020
   "111010010010011010", -- Line 1   Column 421   Coefficient -0.17851257
   "000000001000010100", -- Line 1   Column 422   Coefficient 0.00405884
   "000010001100000001", -- Line 1   Column 423   Coefficient 0.06836700
   "111001011100001110", -- Line 1   Column 424   Coefficient -0.20497131
   "101011001100100000", -- Line 1   Column 425   Coefficient -0.65014648
   "100101100010001110", -- Line 1   Column 426   Coefficient -0.82704163
   "110001001101111000", -- Line 1   Column 427   Coefficient -0.46197510
   "000111101111001000", -- Line 1   Column 428   Coefficient 0.24176025
   "011000100000110011", -- Line 1   Column 429   Coefficient 0.76601410
   "011000010101011011", -- Line 1   Column 430   Coefficient 0.76045990
   "001011010100111000", -- Line 1   Column 431   Coefficient 0.35394287
   "111111100000001001", -- Line 1   Column 432   Coefficient -0.01555634
   "111110001110101111", -- Line 1   Column 433   Coefficient -0.05530548
   "000100000010011110", -- Line 1   Column 434   Coefficient 0.12620544
   "000110101010011000", -- Line 1   Column 435   Coefficient 0.20819092
   "000001100011101000", -- Line 1   Column 436   Coefficient 0.04864502
   "111010100101011001", -- Line 1   Column 437   Coefficient -0.16924286
   "111010000010000111", -- Line 1   Column 438   Coefficient -0.18647003
   "111111101111000001", -- Line 1   Column 439   Coefficient -0.00829315
   "000010010111010110", -- Line 1   Column 440   Coefficient 0.07389832
   "111010010100110101", -- Line 1   Column 441   Coefficient -0.17733002
   "101100000010100100", -- Line 1   Column 442   Coefficient -0.62374878
   "100101011001010011", -- Line 1   Column 443   Coefficient -0.83139801
   "101111111100100011", -- Line 1   Column 444   Coefficient -0.50168610
   "000110001110010001", -- Line 1   Column 445   Coefficient 0.19446564
   "010111110111111000", -- Line 1   Column 446   Coefficient 0.74603271
   "011000110111110111", -- Line 1   Column 447   Coefficient 0.77727509
   "001100010100011100", -- Line 1   Column 448   Coefficient 0.38497925
   "000000000000000000", -- Line 1   Column 449   Coefficient 0.00000000
   "111101111111100010", -- Line 1   Column 450   Coefficient -0.06272888
   "000011101001000111", -- Line 1   Column 451   Coefficient 0.11382294
   "000110101111001111", -- Line 1   Column 452   Coefficient 0.21056366
   "000010000011111010", -- Line 1   Column 453   Coefficient 0.06440735
   "111010111010011110", -- Line 1   Column 454   Coefficient -0.15895081
   "111001110011110110", -- Line 1   Column 455   Coefficient -0.19343567
   "111111010100110011", -- Line 1   Column 456   Coefficient -0.02109528
   "000010011111010100", -- Line 1   Column 457   Coefficient 0.07778931
   "111011001011011000", -- Line 1   Column 458   Coefficient -0.15069580
   "101100111010111010", -- Line 1   Column 459   Coefficient -0.59623718
   "100101010101101100", -- Line 1   Column 460   Coefficient -0.83316040
   "101110101110110111", -- Line 1   Column 461   Coefficient -0.53961945
   "000100101011111110", -- Line 1   Column 462   Coefficient 0.14646912
   "010111001001110011", -- Line 1   Column 463   Coefficient 0.72353363
   "011001010110001010", -- Line 1   Column 464   Coefficient 0.79206848
   "001101010100001011", -- Line 1   Column 465   Coefficient 0.41609955
   "000000100011001001", -- Line 1   Column 466   Coefficient 0.01715851
   "111101110010101110", -- Line 1   Column 467   Coefficient -0.06898499
   "000011001110111000", -- Line 1   Column 468   Coefficient 0.10101318
   "000110110001100100", -- Line 1   Column 469   Coefficient 0.21170044
   "000010100011011000", -- Line 1   Column 470   Coefficient 0.07977295
   "111011010001011111", -- Line 1   Column 471   Coefficient -0.14771271
   "111001100111101111", -- Line 1   Column 472   Coefficient -0.19934845
   "111110111001111010", -- Line 1   Column 473   Coefficient -0.03422546
   "000010100011111110", -- Line 1   Column 474   Coefficient 0.08006287
   "111011111111101011", -- Line 1   Column 475   Coefficient -0.12516022
   "101101110101001111", -- Line 1   Column 476   Coefficient -0.56775665
   "100101010111010100", -- Line 1   Column 477   Coefficient -0.83236694
   "101101100101000100", -- Line 1   Column 478   Coefficient -0.57565308
   "000011001000100101", -- Line 1   Column 479   Coefficient 0.09793854
   "010110010110101011", -- Line 1   Column 480   Coefficient 0.69857025
   "011001110000000111", -- Line 1   Column 481   Coefficient 0.80474091
   "001110010011110010", -- Line 1   Column 482   Coefficient 0.44715881
   "000001001001011111", -- Line 1   Column 483   Coefficient 0.03588104
   "111101101000011110", -- Line 1   Column 484   Coefficient -0.07398987
   "000010110011111110", -- Line 1   Column 485   Coefficient 0.08787537
   "000110110001011010", -- Line 1   Column 486   Coefficient 0.21162415
   "000011000001111000", -- Line 1   Column 487   Coefficient 0.09466553
   "111011101010010100", -- Line 1   Column 488   Coefficient -0.13558960
   "111001011101111001", -- Line 1   Column 489   Coefficient -0.20415497
   "111110011110100011", -- Line 1   Column 490   Coefficient -0.04758453
   "000010100101011011", -- Line 1   Column 491   Coefficient 0.08077240
   "111100110001100001", -- Line 1   Column 492   Coefficient -0.10082245
   "101110110001001111", -- Line 1   Column 493   Coefficient -0.53845978
   "100101011110000100", -- Line 1   Column 494   Coefficient -0.82907104
   "101100011111011001", -- Line 1   Column 495   Coefficient -0.60967255
   "000001100100011110", -- Line 1   Column 496   Coefficient 0.04905701
   "010101011110101011", -- Line 1   Column 497   Coefficient 0.67122650
   "011010000101011111", -- Line 1   Column 498   Coefficient 0.81517792
   "001111010010111101", -- Line 1   Column 499   Coefficient 0.47800446
   "000001110010111010", -- Line 1   Column 500   Coefficient 0.05610657
   "111101100000111011", -- Line 1   Column 501   Coefficient -0.07767487
   "000010011000100111", -- Line 1   Column 502   Coefficient 0.07451630
   "000110101110110000", -- Line 1   Column 503   Coefficient 0.21032715
   "000011011111001110", -- Line 1   Column 504   Coefficient 0.10899353
   "111100000100110011", -- Line 1   Column 505   Coefficient -0.12265778
   "111001010110010111", -- Line 1   Column 506   Coefficient -0.20783234
   "111110000010111110", -- Line 1   Column 507   Coefficient -0.06105042
   "000010100011110000", -- Line 1   Column 508   Coefficient 0.07995605
   "111101100000101101", -- Line 1   Column 509   Coefficient -0.07778168
   "101111101110100111", -- Line 1   Column 510   Coefficient -0.50849152
   "100101101001110110", -- Line 1   Column 511   Coefficient -0.82331848
   "101011011110000110", -- Line 1   Column 512   Coefficient -0.64155579
   "000000000000000000", -- Line 1   Column 513   Coefficient 0.00000000
   "010100100001111010", -- Line 1   Column 514   Coefficient 0.64155579
   "011010010110001010", -- Line 1   Column 515   Coefficient 0.82331848
   "010000010001011001", -- Line 1   Column 516   Coefficient 0.50849152
   "000010011111010011", -- Line 1   Column 517   Coefficient 0.07778168
   "111101011100010000", -- Line 1   Column 518   Coefficient -0.07995605
   "000001111101000010", -- Line 1   Column 519   Coefficient 0.06105042
   "000110101001101001", -- Line 1   Column 520   Coefficient 0.20783234
   "000011111011001101", -- Line 1   Column 521   Coefficient 0.12265778
   "111100100000110010", -- Line 1   Column 522   Coefficient -0.10899353
   "111001010001010000", -- Line 1   Column 523   Coefficient -0.21032715
   "111101100111011001", -- Line 1   Column 524   Coefficient -0.07451630
   "000010011111000101", -- Line 1   Column 525   Coefficient 0.07767487
   "111110001101000110", -- Line 1   Column 526   Coefficient -0.05610657
   "110000101101000011", -- Line 1   Column 527   Coefficient -0.47800446
   "100101111010100001", -- Line 1   Column 528   Coefficient -0.81517792
   "101010100001010101", -- Line 1   Column 529   Coefficient -0.67122650
   "111110011011100010", -- Line 1   Column 530   Coefficient -0.04905701
   "010011100000100111", -- Line 1   Column 531   Coefficient 0.60967255
   "011010100001111100", -- Line 1   Column 532   Coefficient 0.82907104
   "010001001110110001", -- Line 1   Column 533   Coefficient 0.53845978
   "000011001110011111", -- Line 1   Column 534   Coefficient 0.10082245
   "111101011010100101", -- Line 1   Column 535   Coefficient -0.08077240
   "000001100001011101", -- Line 1   Column 536   Coefficient 0.04758453
   "000110100010000111", -- Line 1   Column 537   Coefficient 0.20415497
   "000100010101101100", -- Line 1   Column 538   Coefficient 0.13558960
   "111100111110001000", -- Line 1   Column 539   Coefficient -0.09466553
   "111001001110100110", -- Line 1   Column 540   Coefficient -0.21162415
   "111101001100000010", -- Line 1   Column 541   Coefficient -0.08787537
   "000010010111100010", -- Line 1   Column 542   Coefficient 0.07398987
   "111110110110100001", -- Line 1   Column 543   Coefficient -0.03588104
   "110001101100001110", -- Line 1   Column 544   Coefficient -0.44715881
   "100110001111111001", -- Line 1   Column 545   Coefficient -0.80474091
   "101001101001010101", -- Line 1   Column 546   Coefficient -0.69857025
   "111100110111011011", -- Line 1   Column 547   Coefficient -0.09793854
   "010010011010111100", -- Line 1   Column 548   Coefficient 0.57565308
   "011010101000101100", -- Line 1   Column 549   Coefficient 0.83236694
   "010010001010110001", -- Line 1   Column 550   Coefficient 0.56775665
   "000100000000010101", -- Line 1   Column 551   Coefficient 0.12516022
   "111101011100000010", -- Line 1   Column 552   Coefficient -0.08006287
   "000001000110000110", -- Line 1   Column 553   Coefficient 0.03422546
   "000110011000010001", -- Line 1   Column 554   Coefficient 0.19934845
   "000100101110100001", -- Line 1   Column 555   Coefficient 0.14771271
   "111101011100101000", -- Line 1   Column 556   Coefficient -0.07977295
   "111001001110011100", -- Line 1   Column 557   Coefficient -0.21170044
   "111100110001001000", -- Line 1   Column 558   Coefficient -0.10101318
   "000010001101010010", -- Line 1   Column 559   Coefficient 0.06898499
   "111111011100110111", -- Line 1   Column 560   Coefficient -0.01715851
   "110010101011110101", -- Line 1   Column 561   Coefficient -0.41609955
   "100110101001110110", -- Line 1   Column 562   Coefficient -0.79206848
   "101000110110001101", -- Line 1   Column 563   Coefficient -0.72353363
   "111011010100000010", -- Line 1   Column 564   Coefficient -0.14646912
   "010001010001001001", -- Line 1   Column 565   Coefficient 0.53961945
   "011010101010010100", -- Line 1   Column 566   Coefficient 0.83316040
   "010011000101000110", -- Line 1   Column 567   Coefficient 0.59623718
   "000100110100101000", -- Line 1   Column 568   Coefficient 0.15069580
   "111101100000101100", -- Line 1   Column 569   Coefficient -0.07778931
   "000000101011001101", -- Line 1   Column 570   Coefficient 0.02109528
   "000110001100001010", -- Line 1   Column 571   Coefficient 0.19343567
   "000101000101100010", -- Line 1   Column 572   Coefficient 0.15895081
   "111101111100000110", -- Line 1   Column 573   Coefficient -0.06440735
   "111001010000110001", -- Line 1   Column 574   Coefficient -0.21056366
   "111100010110111001", -- Line 1   Column 575   Coefficient -0.11382294
   "000010000000011110", -- Line 1   Column 576   Coefficient 0.06272888
   "000000000000000000", -- Line 1   Column 577   Coefficient 0.00000000
   "110011101011100100", -- Line 1   Column 578   Coefficient -0.38497925
   "100111001000001001", -- Line 1   Column 579   Coefficient -0.77727509
   "101000001000001000", -- Line 1   Column 580   Coefficient -0.74603271
   "111001110001101111", -- Line 1   Column 581   Coefficient -0.19446564
   "010000000011011101", -- Line 1   Column 582   Coefficient 0.50168610
   "011010100110101101", -- Line 1   Column 583   Coefficient 0.83139801
   "010011111101011100", -- Line 1   Column 584   Coefficient 0.62374878
   "000101101011001011", -- Line 1   Column 585   Coefficient 0.17733002
   "111101101000101010", -- Line 1   Column 586   Coefficient -0.07389832
   "000000010000111111", -- Line 1   Column 587   Coefficient 0.00829315
   "000101111101111001", -- Line 1   Column 588   Coefficient 0.18647003
   "000101011010100111", -- Line 1   Column 589   Coefficient 0.16924286
   "111110011100011000", -- Line 1   Column 590   Coefficient -0.04864502
   "111001010101101000", -- Line 1   Column 591   Coefficient -0.20819092
   "111011111101100010", -- Line 1   Column 592   Coefficient -0.12620544
   "000001110001010001", -- Line 1   Column 593   Coefficient 0.05530548
   "000000011111110111", -- Line 1   Column 594   Coefficient 0.01555634
   "110100101011001000", -- Line 1   Column 595   Coefficient -0.35394287
   "100111101010100101", -- Line 1   Column 596   Coefficient -0.76045990
   "100111011111001101", -- Line 1   Column 597   Coefficient -0.76601410
   "111000010000111000", -- Line 1   Column 598   Coefficient -0.24176025
   "001110110010001000", -- Line 1   Column 599   Coefficient 0.46197510
   "011010011101110010", -- Line 1   Column 600   Coefficient 0.82704163
   "010100110011100000", -- Line 1   Column 601   Coefficient 0.65014648
   "000110100011110010", -- Line 1   Column 602   Coefficient 0.20497131
   "111101110011111111", -- Line 1   Column 603   Coefficient -0.06836700
   "111111110111101100", -- Line 1   Column 604   Coefficient -0.00405884
   "000101101101100110", -- Line 1   Column 605   Coefficient 0.17851257
   "000101101101100111", -- Line 1   Column 606   Coefficient 0.17852020
   "111110111101010000", -- Line 1   Column 607   Coefficient -0.03259277
   "111001011100111110", -- Line 1   Column 608   Coefficient -0.20460510
   "111011100101001111", -- Line 1   Column 609   Coefficient -0.13806915
   "000001011111110111", -- Line 1   Column 610   Coefficient 0.04680634
   "000000111100010110", -- Line 1   Column 611   Coefficient 0.02946472
   "110101101010001101", -- Line 1   Column 612   Coefficient -0.32314301
   "101000010000111100", -- Line 1   Column 613   Coefficient -0.74172974
   "100110111011100001", -- Line 1   Column 614   Coefficient -0.78343964
   "110110110001110010", -- Line 1   Column 615   Coefficient -0.28819275
   "001101011101011101", -- Line 1   Column 616   Coefficient 0.42063141
   "011010001111100001", -- Line 1   Column 617   Coefficient 0.82007599
   "010101100110111110", -- Line 1   Column 618   Coefficient 0.67527771
   "000111011110001100", -- Line 1   Column 619   Coefficient 0.23348999
   "111110000010101111", -- Line 1   Column 620   Coefficient -0.06116486
   "111111011111100010", -- Line 1   Column 621   Coefficient -0.01585388
   "000101011011011000", -- Line 1   Column 622   Coefficient 0.16961670
   "000101111110011101", -- Line 1   Column 623   Coefficient 0.18674469
   "111111011110100001", -- Line 1   Column 624   Coefficient -0.01634979
   "111001100110110001", -- Line 1   Column 625   Coefficient -0.19982147
   "111011001110001101", -- Line 1   Column 626   Coefficient -0.14931488
   "000001001100011101", -- Line 1   Column 627   Coefficient 0.03733063
   "000001010101011100", -- Line 1   Column 628   Coefficient 0.04171753
   "110110101000100010", -- Line 1   Column 629   Coefficient -0.29270935
   "101000111010111110", -- Line 1   Column 630   Coefficient -0.72120667
   "100110011101001001", -- Line 1   Column 631   Coefficient -0.79827118
   "110101010100110101", -- Line 1   Column 632   Coefficient -0.33358002
   "001100000101101101", -- Line 1   Column 633   Coefficient 0.37778473
   "011001111011111000", -- Line 1   Column 634   Coefficient 0.81048584
   "010110010111100101", -- Line 1   Column 635   Coefficient 0.69901276
   "001000011010001011", -- Line 1   Column 636   Coefficient 0.26277924
   "111110010100111011", -- Line 1   Column 637   Coefficient -0.05228424
   "111111001000101111", -- Line 1   Column 638   Coefficient -0.02698517
   "000101000111011001", -- Line 1   Column 639   Coefficient 0.15985870
   "000110001101000001", -- Line 1   Column 640   Coefficient 0.19385529
   "000000000000000000", -- Line 1   Column 641   Coefficient 0.00000000
   "111001110010111111", -- Line 1   Column 642   Coefficient -0.19385529
   "111010111000100111", -- Line 1   Column 643   Coefficient -0.15985870
   "000000110111010001", -- Line 1   Column 644   Coefficient 0.02698517
   "000001101011000101", -- Line 1   Column 645   Coefficient 0.05228424
   "110111100101110101", -- Line 1   Column 646   Coefficient -0.26277924
   "101001101000011011", -- Line 1   Column 647   Coefficient -0.69901276
   "100110000100001000", -- Line 1   Column 648   Coefficient -0.81048584
   "110011111010010011", -- Line 1   Column 649   Coefficient -0.37778473
   "001010101011001011", -- Line 1   Column 650   Coefficient 0.33358002
   "011001100010110111", -- Line 1   Column 651   Coefficient 0.79827118
   "010111000101000010", -- Line 1   Column 652   Coefficient 0.72120667
   "001001010111011110", -- Line 1   Column 653   Coefficient 0.29270935
   "111110101010100100", -- Line 1   Column 654   Coefficient -0.04171753
   "111110110011100011", -- Line 1   Column 655   Coefficient -0.03733063
   "000100110001110011", -- Line 1   Column 656   Coefficient 0.14931488
   "000110011001001111", -- Line 1   Column 657   Coefficient 0.19982147
   "000000100001011111", -- Line 1   Column 658   Coefficient 0.01634979
   "111010000001100011", -- Line 1   Column 659   Coefficient -0.18674469
   "111010100100101000", -- Line 1   Column 660   Coefficient -0.16961670
   "000000100000011110", -- Line 1   Column 661   Coefficient 0.01585388
   "000001111101010001", -- Line 1   Column 662   Coefficient 0.06116486
   "111000100001110100", -- Line 1   Column 663   Coefficient -0.23348999
   "101010011001000010", -- Line 1   Column 664   Coefficient -0.67527771
   "100101110000011111", -- Line 1   Column 665   Coefficient -0.82007599
   "110010100010100011", -- Line 1   Column 666   Coefficient -0.42063141
   "001001001110001110", -- Line 1   Column 667   Coefficient 0.28819275
   "011001000100011111", -- Line 1   Column 668   Coefficient 0.78343964
   "010111101111000100", -- Line 1   Column 669   Coefficient 0.74172974
   "001010010101110011", -- Line 1   Column 670   Coefficient 0.32314301
   "111111000011101010", -- Line 1   Column 671   Coefficient -0.02946472
   "111110100000001001", -- Line 1   Column 672   Coefficient -0.04680634
   "000100011010110001", -- Line 1   Column 673   Coefficient 0.13806915
   "000110100011000010", -- Line 1   Column 674   Coefficient 0.20460510
   "000001000010110000", -- Line 1   Column 675   Coefficient 0.03259277
   "111010010010011001", -- Line 1   Column 676   Coefficient -0.17852020
   "111010010010011010", -- Line 1   Column 677   Coefficient -0.17851257
   "000000001000010100", -- Line 1   Column 678   Coefficient 0.00405884
   "000010001100000001", -- Line 1   Column 679   Coefficient 0.06836700
   "111001011100001110", -- Line 1   Column 680   Coefficient -0.20497131
   "101011001100100000", -- Line 1   Column 681   Coefficient -0.65014648
   "100101100010001110", -- Line 1   Column 682   Coefficient -0.82704163
   "110001001101111000", -- Line 1   Column 683   Coefficient -0.46197510
   "000111101111001000", -- Line 1   Column 684   Coefficient 0.24176025
   "011000100000110011", -- Line 1   Column 685   Coefficient 0.76601410
   "011000010101011011", -- Line 1   Column 686   Coefficient 0.76045990
   "001011010100111000", -- Line 1   Column 687   Coefficient 0.35394287
   "111111100000001001", -- Line 1   Column 688   Coefficient -0.01555634
   "111110001110101111", -- Line 1   Column 689   Coefficient -0.05530548
   "000100000010011110", -- Line 1   Column 690   Coefficient 0.12620544
   "000110101010011000", -- Line 1   Column 691   Coefficient 0.20819092
   "000001100011101000", -- Line 1   Column 692   Coefficient 0.04864502
   "111010100101011001", -- Line 1   Column 693   Coefficient -0.16924286
   "111010000010000111", -- Line 1   Column 694   Coefficient -0.18647003
   "111111101111000001", -- Line 1   Column 695   Coefficient -0.00829315
   "000010010111010110", -- Line 1   Column 696   Coefficient 0.07389832
   "111010010100110101", -- Line 1   Column 697   Coefficient -0.17733002
   "101100000010100100", -- Line 1   Column 698   Coefficient -0.62374878
   "100101011001010011", -- Line 1   Column 699   Coefficient -0.83139801
   "101111111100100011", -- Line 1   Column 700   Coefficient -0.50168610
   "000110001110010001", -- Line 1   Column 701   Coefficient 0.19446564
   "010111110111111000", -- Line 1   Column 702   Coefficient 0.74603271
   "011000110111110111", -- Line 1   Column 703   Coefficient 0.77727509
   "001100010100011100", -- Line 1   Column 704   Coefficient 0.38497925
   "000000000000000000", -- Line 1   Column 705   Coefficient 0.00000000
   "111101111111100010", -- Line 1   Column 706   Coefficient -0.06272888
   "000011101001000111", -- Line 1   Column 707   Coefficient 0.11382294
   "000110101111001111", -- Line 1   Column 708   Coefficient 0.21056366
   "000010000011111010", -- Line 1   Column 709   Coefficient 0.06440735
   "111010111010011110", -- Line 1   Column 710   Coefficient -0.15895081
   "111001110011110110", -- Line 1   Column 711   Coefficient -0.19343567
   "111111010100110011", -- Line 1   Column 712   Coefficient -0.02109528
   "000010011111010100", -- Line 1   Column 713   Coefficient 0.07778931
   "111011001011011000", -- Line 1   Column 714   Coefficient -0.15069580
   "101100111010111010", -- Line 1   Column 715   Coefficient -0.59623718
   "100101010101101100", -- Line 1   Column 716   Coefficient -0.83316040
   "101110101110110111", -- Line 1   Column 717   Coefficient -0.53961945
   "000100101011111110", -- Line 1   Column 718   Coefficient 0.14646912
   "010111001001110011", -- Line 1   Column 719   Coefficient 0.72353363
   "011001010110001010", -- Line 1   Column 720   Coefficient 0.79206848
   "001101010100001011", -- Line 1   Column 721   Coefficient 0.41609955
   "000000100011001001", -- Line 1   Column 722   Coefficient 0.01715851
   "111101110010101110", -- Line 1   Column 723   Coefficient -0.06898499
   "000011001110111000", -- Line 1   Column 724   Coefficient 0.10101318
   "000110110001100100", -- Line 1   Column 725   Coefficient 0.21170044
   "000010100011011000", -- Line 1   Column 726   Coefficient 0.07977295
   "111011010001011111", -- Line 1   Column 727   Coefficient -0.14771271
   "111001100111101111", -- Line 1   Column 728   Coefficient -0.19934845
   "111110111001111010", -- Line 1   Column 729   Coefficient -0.03422546
   "000010100011111110", -- Line 1   Column 730   Coefficient 0.08006287
   "111011111111101011", -- Line 1   Column 731   Coefficient -0.12516022
   "101101110101001111", -- Line 1   Column 732   Coefficient -0.56775665
   "100101010111010100", -- Line 1   Column 733   Coefficient -0.83236694
   "101101100101000100", -- Line 1   Column 734   Coefficient -0.57565308
   "000011001000100101", -- Line 1   Column 735   Coefficient 0.09793854
   "010110010110101011", -- Line 1   Column 736   Coefficient 0.69857025
   "011001110000000111", -- Line 1   Column 737   Coefficient 0.80474091
   "001110010011110010", -- Line 1   Column 738   Coefficient 0.44715881
   "000001001001011111", -- Line 1   Column 739   Coefficient 0.03588104
   "111101101000011110", -- Line 1   Column 740   Coefficient -0.07398987
   "000010110011111110", -- Line 1   Column 741   Coefficient 0.08787537
   "000110110001011010", -- Line 1   Column 742   Coefficient 0.21162415
   "000011000001111000", -- Line 1   Column 743   Coefficient 0.09466553
   "111011101010010100", -- Line 1   Column 744   Coefficient -0.13558960
   "111001011101111001", -- Line 1   Column 745   Coefficient -0.20415497
   "111110011110100011", -- Line 1   Column 746   Coefficient -0.04758453
   "000010100101011011", -- Line 1   Column 747   Coefficient 0.08077240
   "111100110001100001", -- Line 1   Column 748   Coefficient -0.10082245
   "101110110001001111", -- Line 1   Column 749   Coefficient -0.53845978
   "100101011110000100", -- Line 1   Column 750   Coefficient -0.82907104
   "101100011111011001", -- Line 1   Column 751   Coefficient -0.60967255
   "000001100100011110", -- Line 1   Column 752   Coefficient 0.04905701
   "010101011110101011", -- Line 1   Column 753   Coefficient 0.67122650
   "011010000101011111", -- Line 1   Column 754   Coefficient 0.81517792
   "001111010010111101", -- Line 1   Column 755   Coefficient 0.47800446
   "000001110010111010", -- Line 1   Column 756   Coefficient 0.05610657
   "111101100000111011", -- Line 1   Column 757   Coefficient -0.07767487
   "000010011000100111", -- Line 1   Column 758   Coefficient 0.07451630
   "000110101110110000", -- Line 1   Column 759   Coefficient 0.21032715
   "000011011111001110", -- Line 1   Column 760   Coefficient 0.10899353
   "111100000100110011", -- Line 1   Column 761   Coefficient -0.12265778
   "111001010110010111", -- Line 1   Column 762   Coefficient -0.20783234
   "111110000010111110", -- Line 1   Column 763   Coefficient -0.06105042
   "000010100011110000", -- Line 1   Column 764   Coefficient 0.07995605
   "111101100000101101", -- Line 1   Column 765   Coefficient -0.07778168
   "101111101110100111", -- Line 1   Column 766   Coefficient -0.50849152
   "100101101001110110", -- Line 1   Column 767   Coefficient -0.82331848
   "101011011110000110", -- Line 1   Column 768   Coefficient -0.64155579
   "000000000000000000", -- Line 1   Column 769   Coefficient 0.00000000
   "010100100001111010", -- Line 1   Column 770   Coefficient 0.64155579
   "011010010110001010", -- Line 1   Column 771   Coefficient 0.82331848
   "010000010001011001", -- Line 1   Column 772   Coefficient 0.50849152
   "000010011111010011", -- Line 1   Column 773   Coefficient 0.07778168
   "111101011100010000", -- Line 1   Column 774   Coefficient -0.07995605
   "000001111101000010", -- Line 1   Column 775   Coefficient 0.06105042
   "000110101001101001", -- Line 1   Column 776   Coefficient 0.20783234
   "000011111011001101", -- Line 1   Column 777   Coefficient 0.12265778
   "111100100000110010", -- Line 1   Column 778   Coefficient -0.10899353
   "111001010001010000", -- Line 1   Column 779   Coefficient -0.21032715
   "111101100111011001", -- Line 1   Column 780   Coefficient -0.07451630
   "000010011111000101", -- Line 1   Column 781   Coefficient 0.07767487
   "111110001101000110", -- Line 1   Column 782   Coefficient -0.05610657
   "110000101101000011", -- Line 1   Column 783   Coefficient -0.47800446
   "100101111010100001", -- Line 1   Column 784   Coefficient -0.81517792
   "101010100001010101", -- Line 1   Column 785   Coefficient -0.67122650
   "111110011011100010", -- Line 1   Column 786   Coefficient -0.04905701
   "010011100000100111", -- Line 1   Column 787   Coefficient 0.60967255
   "011010100001111100", -- Line 1   Column 788   Coefficient 0.82907104
   "010001001110110001", -- Line 1   Column 789   Coefficient 0.53845978
   "000011001110011111", -- Line 1   Column 790   Coefficient 0.10082245
   "111101011010100101", -- Line 1   Column 791   Coefficient -0.08077240
   "000001100001011101", -- Line 1   Column 792   Coefficient 0.04758453
   "000110100010000111", -- Line 1   Column 793   Coefficient 0.20415497
   "000100010101101100", -- Line 1   Column 794   Coefficient 0.13558960
   "111100111110001000", -- Line 1   Column 795   Coefficient -0.09466553
   "111001001110100110", -- Line 1   Column 796   Coefficient -0.21162415
   "111101001100000010", -- Line 1   Column 797   Coefficient -0.08787537
   "000010010111100010", -- Line 1   Column 798   Coefficient 0.07398987
   "111110110110100001", -- Line 1   Column 799   Coefficient -0.03588104
   "110001101100001110", -- Line 1   Column 800   Coefficient -0.44715881
   "100110001111111001", -- Line 1   Column 801   Coefficient -0.80474091
   "101001101001010101", -- Line 1   Column 802   Coefficient -0.69857025
   "111100110111011011", -- Line 1   Column 803   Coefficient -0.09793854
   "010010011010111100", -- Line 1   Column 804   Coefficient 0.57565308
   "011010101000101100", -- Line 1   Column 805   Coefficient 0.83236694
   "010010001010110001", -- Line 1   Column 806   Coefficient 0.56775665
   "000100000000010101", -- Line 1   Column 807   Coefficient 0.12516022
   "111101011100000010", -- Line 1   Column 808   Coefficient -0.08006287
   "000001000110000110", -- Line 1   Column 809   Coefficient 0.03422546
   "000110011000010001", -- Line 1   Column 810   Coefficient 0.19934845
   "000100101110100001", -- Line 1   Column 811   Coefficient 0.14771271
   "111101011100101000", -- Line 1   Column 812   Coefficient -0.07977295
   "111001001110011100", -- Line 1   Column 813   Coefficient -0.21170044
   "111100110001001000", -- Line 1   Column 814   Coefficient -0.10101318
   "000010001101010010", -- Line 1   Column 815   Coefficient 0.06898499
   "111111011100110111", -- Line 1   Column 816   Coefficient -0.01715851
   "110010101011110101", -- Line 1   Column 817   Coefficient -0.41609955
   "100110101001110110", -- Line 1   Column 818   Coefficient -0.79206848
   "101000110110001101", -- Line 1   Column 819   Coefficient -0.72353363
   "111011010100000010", -- Line 1   Column 820   Coefficient -0.14646912
   "010001010001001001", -- Line 1   Column 821   Coefficient 0.53961945
   "011010101010010100", -- Line 1   Column 822   Coefficient 0.83316040
   "010011000101000110", -- Line 1   Column 823   Coefficient 0.59623718
   "000100110100101000", -- Line 1   Column 824   Coefficient 0.15069580
   "111101100000101100", -- Line 1   Column 825   Coefficient -0.07778931
   "000000101011001101", -- Line 1   Column 826   Coefficient 0.02109528
   "000110001100001010", -- Line 1   Column 827   Coefficient 0.19343567
   "000101000101100010", -- Line 1   Column 828   Coefficient 0.15895081
   "111101111100000110", -- Line 1   Column 829   Coefficient -0.06440735
   "111001010000110001", -- Line 1   Column 830   Coefficient -0.21056366
   "111100010110111001", -- Line 1   Column 831   Coefficient -0.11382294
   "000010000000011110", -- Line 1   Column 832   Coefficient 0.06272888
   "000000000000000000", -- Line 1   Column 833   Coefficient 0.00000000
   "110011101011100100", -- Line 1   Column 834   Coefficient -0.38497925
   "100111001000001001", -- Line 1   Column 835   Coefficient -0.77727509
   "101000001000001000", -- Line 1   Column 836   Coefficient -0.74603271
   "111001110001101111", -- Line 1   Column 837   Coefficient -0.19446564
   "010000000011011101", -- Line 1   Column 838   Coefficient 0.50168610
   "011010100110101101", -- Line 1   Column 839   Coefficient 0.83139801
   "010011111101011100", -- Line 1   Column 840   Coefficient 0.62374878
   "000101101011001011", -- Line 1   Column 841   Coefficient 0.17733002
   "111101101000101010", -- Line 1   Column 842   Coefficient -0.07389832
   "000000010000111111", -- Line 1   Column 843   Coefficient 0.00829315
   "000101111101111001", -- Line 1   Column 844   Coefficient 0.18647003
   "000101011010100111", -- Line 1   Column 845   Coefficient 0.16924286
   "111110011100011000", -- Line 1   Column 846   Coefficient -0.04864502
   "111001010101101000", -- Line 1   Column 847   Coefficient -0.20819092
   "111011111101100010", -- Line 1   Column 848   Coefficient -0.12620544
   "000001110001010001", -- Line 1   Column 849   Coefficient 0.05530548
   "000000011111110111", -- Line 1   Column 850   Coefficient 0.01555634
   "110100101011001000", -- Line 1   Column 851   Coefficient -0.35394287
   "100111101010100101", -- Line 1   Column 852   Coefficient -0.76045990
   "100111011111001101", -- Line 1   Column 853   Coefficient -0.76601410
   "111000010000111000", -- Line 1   Column 854   Coefficient -0.24176025
   "001110110010001000", -- Line 1   Column 855   Coefficient 0.46197510
   "011010011101110010", -- Line 1   Column 856   Coefficient 0.82704163
   "010100110011100000", -- Line 1   Column 857   Coefficient 0.65014648
   "000110100011110010", -- Line 1   Column 858   Coefficient 0.20497131
   "111101110011111111", -- Line 1   Column 859   Coefficient -0.06836700
   "111111110111101100", -- Line 1   Column 860   Coefficient -0.00405884
   "000101101101100110", -- Line 1   Column 861   Coefficient 0.17851257
   "000101101101100111", -- Line 1   Column 862   Coefficient 0.17852020
   "111110111101010000", -- Line 1   Column 863   Coefficient -0.03259277
   "111001011100111110", -- Line 1   Column 864   Coefficient -0.20460510
   "111011100101001111", -- Line 1   Column 865   Coefficient -0.13806915
   "000001011111110111", -- Line 1   Column 866   Coefficient 0.04680634
   "000000111100010110", -- Line 1   Column 867   Coefficient 0.02946472
   "110101101010001101", -- Line 1   Column 868   Coefficient -0.32314301
   "101000010000111100", -- Line 1   Column 869   Coefficient -0.74172974
   "100110111011100001", -- Line 1   Column 870   Coefficient -0.78343964
   "110110110001110010", -- Line 1   Column 871   Coefficient -0.28819275
   "001101011101011101", -- Line 1   Column 872   Coefficient 0.42063141
   "011010001111100001", -- Line 1   Column 873   Coefficient 0.82007599
   "010101100110111110", -- Line 1   Column 874   Coefficient 0.67527771
   "000111011110001100", -- Line 1   Column 875   Coefficient 0.23348999
   "111110000010101111", -- Line 1   Column 876   Coefficient -0.06116486
   "111111011111100010", -- Line 1   Column 877   Coefficient -0.01585388
   "000101011011011000", -- Line 1   Column 878   Coefficient 0.16961670
   "000101111110011101", -- Line 1   Column 879   Coefficient 0.18674469
   "111111011110100001", -- Line 1   Column 880   Coefficient -0.01634979
   "111001100110110001", -- Line 1   Column 881   Coefficient -0.19982147
   "111011001110001101", -- Line 1   Column 882   Coefficient -0.14931488
   "000001001100011101", -- Line 1   Column 883   Coefficient 0.03733063
   "000001010101011100", -- Line 1   Column 884   Coefficient 0.04171753
   "110110101000100010", -- Line 1   Column 885   Coefficient -0.29270935
   "101000111010111110", -- Line 1   Column 886   Coefficient -0.72120667
   "100110011101001001", -- Line 1   Column 887   Coefficient -0.79827118
   "110101010100110101", -- Line 1   Column 888   Coefficient -0.33358002
   "001100000101101101", -- Line 1   Column 889   Coefficient 0.37778473
   "011001111011111000", -- Line 1   Column 890   Coefficient 0.81048584
   "010110010111100101", -- Line 1   Column 891   Coefficient 0.69901276
   "001000011010001011", -- Line 1   Column 892   Coefficient 0.26277924
   "111110010100111011", -- Line 1   Column 893   Coefficient -0.05228424
   "111111001000101111", -- Line 1   Column 894   Coefficient -0.02698517
   "000101000111011001", -- Line 1   Column 895   Coefficient 0.15985870
   "000110001101000001", -- Line 1   Column 896   Coefficient 0.19385529
   "000000000000000000", -- Line 1   Column 897   Coefficient 0.00000000
   "111001110010111111", -- Line 1   Column 898   Coefficient -0.19385529
   "111010111000100111", -- Line 1   Column 899   Coefficient -0.15985870
   "000000110111010001", -- Line 1   Column 900   Coefficient 0.02698517
   "000001101011000101", -- Line 1   Column 901   Coefficient 0.05228424
   "110111100101110101", -- Line 1   Column 902   Coefficient -0.26277924
   "101001101000011011", -- Line 1   Column 903   Coefficient -0.69901276
   "100110000100001000", -- Line 1   Column 904   Coefficient -0.81048584
   "110011111010010011", -- Line 1   Column 905   Coefficient -0.37778473
   "001010101011001011", -- Line 1   Column 906   Coefficient 0.33358002
   "011001100010110111", -- Line 1   Column 907   Coefficient 0.79827118
   "010111000101000010", -- Line 1   Column 908   Coefficient 0.72120667
   "001001010111011110", -- Line 1   Column 909   Coefficient 0.29270935
   "111110101010100100", -- Line 1   Column 910   Coefficient -0.04171753
   "111110110011100011", -- Line 1   Column 911   Coefficient -0.03733063
   "000100110001110011", -- Line 1   Column 912   Coefficient 0.14931488
   "000110011001001111", -- Line 1   Column 913   Coefficient 0.19982147
   "000000100001011111", -- Line 1   Column 914   Coefficient 0.01634979
   "111010000001100011", -- Line 1   Column 915   Coefficient -0.18674469
   "111010100100101000", -- Line 1   Column 916   Coefficient -0.16961670
   "000000100000011110", -- Line 1   Column 917   Coefficient 0.01585388
   "000001111101010001", -- Line 1   Column 918   Coefficient 0.06116486
   "111000100001110100", -- Line 1   Column 919   Coefficient -0.23348999
   "101010011001000010", -- Line 1   Column 920   Coefficient -0.67527771
   "100101110000011111", -- Line 1   Column 921   Coefficient -0.82007599
   "110010100010100011", -- Line 1   Column 922   Coefficient -0.42063141
   "001001001110001110", -- Line 1   Column 923   Coefficient 0.28819275
   "011001000100011111", -- Line 1   Column 924   Coefficient 0.78343964
   "010111101111000100", -- Line 1   Column 925   Coefficient 0.74172974
   "001010010101110011", -- Line 1   Column 926   Coefficient 0.32314301
   "111111000011101010", -- Line 1   Column 927   Coefficient -0.02946472
   "111110100000001001", -- Line 1   Column 928   Coefficient -0.04680634
   "000100011010110001", -- Line 1   Column 929   Coefficient 0.13806915
   "000110100011000010", -- Line 1   Column 930   Coefficient 0.20460510
   "000001000010110000", -- Line 1   Column 931   Coefficient 0.03259277
   "111010010010011001", -- Line 1   Column 932   Coefficient -0.17852020
   "111010010010011010", -- Line 1   Column 933   Coefficient -0.17851257
   "000000001000010100", -- Line 1   Column 934   Coefficient 0.00405884
   "000010001100000001", -- Line 1   Column 935   Coefficient 0.06836700
   "111001011100001110", -- Line 1   Column 936   Coefficient -0.20497131
   "101011001100100000", -- Line 1   Column 937   Coefficient -0.65014648
   "100101100010001110", -- Line 1   Column 938   Coefficient -0.82704163
   "110001001101111000", -- Line 1   Column 939   Coefficient -0.46197510
   "000111101111001000", -- Line 1   Column 940   Coefficient 0.24176025
   "011000100000110011", -- Line 1   Column 941   Coefficient 0.76601410
   "011000010101011011", -- Line 1   Column 942   Coefficient 0.76045990
   "001011010100111000", -- Line 1   Column 943   Coefficient 0.35394287
   "111111100000001001", -- Line 1   Column 944   Coefficient -0.01555634
   "111110001110101111", -- Line 1   Column 945   Coefficient -0.05530548
   "000100000010011110", -- Line 1   Column 946   Coefficient 0.12620544
   "000110101010011000", -- Line 1   Column 947   Coefficient 0.20819092
   "000001100011101000", -- Line 1   Column 948   Coefficient 0.04864502
   "111010100101011001", -- Line 1   Column 949   Coefficient -0.16924286
   "111010000010000111", -- Line 1   Column 950   Coefficient -0.18647003
   "111111101111000001", -- Line 1   Column 951   Coefficient -0.00829315
   "000010010111010110", -- Line 1   Column 952   Coefficient 0.07389832
   "111010010100110101", -- Line 1   Column 953   Coefficient -0.17733002
   "101100000010100100", -- Line 1   Column 954   Coefficient -0.62374878
   "100101011001010011", -- Line 1   Column 955   Coefficient -0.83139801
   "101111111100100011", -- Line 1   Column 956   Coefficient -0.50168610
   "000110001110010001", -- Line 1   Column 957   Coefficient 0.19446564
   "010111110111111000", -- Line 1   Column 958   Coefficient 0.74603271
   "011000110111110111", -- Line 1   Column 959   Coefficient 0.77727509
   "001100010100011100", -- Line 1   Column 960   Coefficient 0.38497925
   "000000000000000000", -- Line 1   Column 961   Coefficient 0.00000000
   "111101111111100010", -- Line 1   Column 962   Coefficient -0.06272888
   "000011101001000111", -- Line 1   Column 963   Coefficient 0.11382294
   "000110101111001111", -- Line 1   Column 964   Coefficient 0.21056366
   "000010000011111010", -- Line 1   Column 965   Coefficient 0.06440735
   "111010111010011110", -- Line 1   Column 966   Coefficient -0.15895081
   "111001110011110110", -- Line 1   Column 967   Coefficient -0.19343567
   "111111010100110011", -- Line 1   Column 968   Coefficient -0.02109528
   "000010011111010100", -- Line 1   Column 969   Coefficient 0.07778931
   "111011001011011000", -- Line 1   Column 970   Coefficient -0.15069580
   "101100111010111010", -- Line 1   Column 971   Coefficient -0.59623718
   "100101010101101100", -- Line 1   Column 972   Coefficient -0.83316040
   "101110101110110111", -- Line 1   Column 973   Coefficient -0.53961945
   "000100101011111110", -- Line 1   Column 974   Coefficient 0.14646912
   "010111001001110011", -- Line 1   Column 975   Coefficient 0.72353363
   "011001010110001010", -- Line 1   Column 976   Coefficient 0.79206848
   "001101010100001011", -- Line 1   Column 977   Coefficient 0.41609955
   "000000100011001001", -- Line 1   Column 978   Coefficient 0.01715851
   "111101110010101110", -- Line 1   Column 979   Coefficient -0.06898499
   "000011001110111000", -- Line 1   Column 980   Coefficient 0.10101318
   "000110110001100100", -- Line 1   Column 981   Coefficient 0.21170044
   "000010100011011000", -- Line 1   Column 982   Coefficient 0.07977295
   "111011010001011111", -- Line 1   Column 983   Coefficient -0.14771271
   "111001100111101111", -- Line 1   Column 984   Coefficient -0.19934845
   "111110111001111010", -- Line 1   Column 985   Coefficient -0.03422546
   "000010100011111110", -- Line 1   Column 986   Coefficient 0.08006287
   "111011111111101011", -- Line 1   Column 987   Coefficient -0.12516022
   "101101110101001111", -- Line 1   Column 988   Coefficient -0.56775665
   "100101010111010100", -- Line 1   Column 989   Coefficient -0.83236694
   "101101100101000100", -- Line 1   Column 990   Coefficient -0.57565308
   "000011001000100101", -- Line 1   Column 991   Coefficient 0.09793854
   "010110010110101011", -- Line 1   Column 992   Coefficient 0.69857025
   "011001110000000111", -- Line 1   Column 993   Coefficient 0.80474091
   "001110010011110010", -- Line 1   Column 994   Coefficient 0.44715881
   "000001001001011111", -- Line 1   Column 995   Coefficient 0.03588104
   "111101101000011110", -- Line 1   Column 996   Coefficient -0.07398987
   "000010110011111110", -- Line 1   Column 997   Coefficient 0.08787537
   "000110110001011010", -- Line 1   Column 998   Coefficient 0.21162415
   "000011000001111000", -- Line 1   Column 999   Coefficient 0.09466553
   "111011101010010100", -- Line 1   Column 1000   Coefficient -0.13558960
   "111001011101111001", -- Line 1   Column 1001   Coefficient -0.20415497
   "111110011110100011", -- Line 1   Column 1002   Coefficient -0.04758453
   "000010100101011011", -- Line 1   Column 1003   Coefficient 0.08077240
   "111100110001100001", -- Line 1   Column 1004   Coefficient -0.10082245
   "101110110001001111", -- Line 1   Column 1005   Coefficient -0.53845978
   "100101011110000100", -- Line 1   Column 1006   Coefficient -0.82907104
   "101100011111011001", -- Line 1   Column 1007   Coefficient -0.60967255
   "000001100100011110", -- Line 1   Column 1008   Coefficient 0.04905701
   "010101011110101011", -- Line 1   Column 1009   Coefficient 0.67122650
   "011010000101011111", -- Line 1   Column 1010   Coefficient 0.81517792
   "001111010010111101", -- Line 1   Column 1011   Coefficient 0.47800446
   "000001110010111010", -- Line 1   Column 1012   Coefficient 0.05610657
   "111101100000111011", -- Line 1   Column 1013   Coefficient -0.07767487
   "000010011000100111", -- Line 1   Column 1014   Coefficient 0.07451630
   "000110101110110000", -- Line 1   Column 1015   Coefficient 0.21032715
   "000011011111001110", -- Line 1   Column 1016   Coefficient 0.10899353
   "111100000100110011", -- Line 1   Column 1017   Coefficient -0.12265778
   "111001010110010111", -- Line 1   Column 1018   Coefficient -0.20783234
   "111110000010111110", -- Line 1   Column 1019   Coefficient -0.06105042
   "000010100011110000", -- Line 1   Column 1020   Coefficient 0.07995605
   "111101100000101101", -- Line 1   Column 1021   Coefficient -0.07778168
   "101111101110100111", -- Line 1   Column 1022   Coefficient -0.50849152
   "100101101001110110", -- Line 1   Column 1023   Coefficient -0.82331848
   "101011011110000110" -- Line 1   Column 1024   Coefficient -0.64155579
);
begin
	process(clk)
	begin
	if(rising_edge(CLK)) then
		A <= rom(to_integer(unsigned(I)));
	end if;
	end process;
end ROM;
