-- IDWT matrix coefficients
--
-- FI - UAQ
--
-- Electronica Avanzada III
--
-- Rene Romero Troncoso
--

library IEEE;
use IEEE.std_logic_1164.all;

entity ROM_IDWT is
   port(
      I : in  std_logic_vector(11 downto 0);
      A : out std_logic_vector(17 downto 0)
      );
   end ROM_IDWT;

architecture LUTable of ROM_IDWT is
begin
   process(I)
   begin
      case I is
         -- Coefficient format 0.18
         when "000000000000" => A <= "000000000000000000"; -- Line 1   Column 1   Coefficient 0.00000000
         when "000000000001" => A <= "000000000000000000"; -- Line 1   Column 2   Coefficient 0.00000000
         when "000000000010" => A <= "000000000000000000"; -- Line 1   Column 3   Coefficient 0.00000000
         when "000000000011" => A <= "000000000000000000"; -- Line 1   Column 4   Coefficient 0.00000000
         when "000000000100" => A <= "000000000000000000"; -- Line 1   Column 5   Coefficient 0.00000000
         when "000000000101" => A <= "000000000000000000"; -- Line 1   Column 6   Coefficient 0.00000000
         when "000000000110" => A <= "000000000000000000"; -- Line 1   Column 7   Coefficient 0.00000000
         when "000000000111" => A <= "000000000000000000"; -- Line 1   Column 8   Coefficient 0.00000000
         when "000000001000" => A <= "000000000000000000"; -- Line 1   Column 9   Coefficient 0.00000000
         when "000000001001" => A <= "000000000000000000"; -- Line 1   Column 10   Coefficient 0.00000000
         when "000000001010" => A <= "000000001101001100"; -- Line 1   Column 11   Coefficient 0.00321960
         when "000000001011" => A <= "111101100010001110"; -- Line 1   Column 12   Coefficient -0.03852081
         when "000000001100" => A <= "010000111010100101"; -- Line 1   Column 13   Coefficient 0.26430130
         when "000000001101" => A <= "000000111110100110"; -- Line 1   Column 14   Coefficient 0.01528168
         when "000000001110" => A <= "000000010110010000"; -- Line 1   Column 15   Coefficient 0.00543213
         when "000000001111" => A <= "000000000001001011"; -- Line 1   Column 16   Coefficient 0.00028610
         when "000000010000" => A <= "000000000000000000"; -- Line 2   Column 1   Coefficient 0.00000000
         when "000000010001" => A <= "000000000000000000"; -- Line 2   Column 2   Coefficient 0.00000000
         when "000000010010" => A <= "000000000000000000"; -- Line 2   Column 3   Coefficient 0.00000000
         when "000000010011" => A <= "000000000000000000"; -- Line 2   Column 4   Coefficient 0.00000000
         when "000000010100" => A <= "000000000000000000"; -- Line 2   Column 5   Coefficient 0.00000000
         when "000000010101" => A <= "000000000000000000"; -- Line 2   Column 6   Coefficient 0.00000000
         when "000000010110" => A <= "000000000000000000"; -- Line 2   Column 7   Coefficient 0.00000000
         when "000000010111" => A <= "000000000000000000"; -- Line 2   Column 8   Coefficient 0.00000000
         when "000000011000" => A <= "000000000000000000"; -- Line 2   Column 9   Coefficient 0.00000000
         when "000000011001" => A <= "000000000000000000"; -- Line 2   Column 10   Coefficient 0.00000000
         when "000000011010" => A <= "000000001010110110"; -- Line 2   Column 11   Coefficient 0.00264740
         when "000000011011" => A <= "111101100010101111"; -- Line 2   Column 12   Coefficient -0.03839493
         when "000000011100" => A <= "001111111010100001"; -- Line 2   Column 13   Coefficient 0.24866104
         when "000000011101" => A <= "000010000100001011"; -- Line 2   Column 14   Coefficient 0.03226852
         when "000000011110" => A <= "000000010100110111"; -- Line 2   Column 15   Coefficient 0.00509262
         when "000000011111" => A <= "111111111110110111"; -- Line 2   Column 16   Coefficient -0.00027847
         when "000000100000" => A <= "111111111111111111"; -- Line 3   Column 1   Coefficient -0.00000381
         when "000000100001" => A <= "000000000000000000"; -- Line 3   Column 2   Coefficient 0.00000000
         when "000000100010" => A <= "000000000000000000"; -- Line 3   Column 3   Coefficient 0.00000000
         when "000000100011" => A <= "000000000000000000"; -- Line 3   Column 4   Coefficient 0.00000000
         when "000000100100" => A <= "000000000000000000"; -- Line 3   Column 5   Coefficient 0.00000000
         when "000000100101" => A <= "000000000000000000"; -- Line 3   Column 6   Coefficient 0.00000000
         when "000000100110" => A <= "000000000000000000"; -- Line 3   Column 7   Coefficient 0.00000000
         when "000000100111" => A <= "000000000000000000"; -- Line 3   Column 8   Coefficient 0.00000000
         when "000000101000" => A <= "000000000000000000"; -- Line 3   Column 9   Coefficient 0.00000000
         when "000000101001" => A <= "000000000000000000"; -- Line 3   Column 10   Coefficient 0.00000000
         when "000000101010" => A <= "000000001000010011"; -- Line 3   Column 11   Coefficient 0.00202560
         when "000000101011" => A <= "111101100110110000"; -- Line 3   Column 12   Coefficient -0.03741455
         when "000000101100" => A <= "001110110101010100"; -- Line 3   Column 13   Coefficient 0.23176575
         when "000000101101" => A <= "000011001010010011"; -- Line 3   Column 14   Coefficient 0.04938889
         when "000000101110" => A <= "000000010100111001"; -- Line 3   Column 15   Coefficient 0.00510025
         when "000000101111" => A <= "111111111100011110"; -- Line 3   Column 16   Coefficient -0.00086212
         when "000000110000" => A <= "000000000000000011"; -- Line 4   Column 1   Coefficient 0.00001144
         when "000000110001" => A <= "000000000000000000"; -- Line 4   Column 2   Coefficient 0.00000000
         when "000000110010" => A <= "000000000000000000"; -- Line 4   Column 3   Coefficient 0.00000000
         when "000000110011" => A <= "000000000000000000"; -- Line 4   Column 4   Coefficient 0.00000000
         when "000000110100" => A <= "000000000000000000"; -- Line 4   Column 5   Coefficient 0.00000000
         when "000000110101" => A <= "000000000000000000"; -- Line 4   Column 6   Coefficient 0.00000000
         when "000000110110" => A <= "000000000000000000"; -- Line 4   Column 7   Coefficient 0.00000000
         when "000000110111" => A <= "000000000000000000"; -- Line 4   Column 8   Coefficient 0.00000000
         when "000000111000" => A <= "000000000000000000"; -- Line 4   Column 9   Coefficient 0.00000000
         when "000000111001" => A <= "000000000000000000"; -- Line 4   Column 10   Coefficient 0.00000000
         when "000000111010" => A <= "000000000011111000"; -- Line 4   Column 11   Coefficient 0.00094604
         when "000000111011" => A <= "111101110100001010"; -- Line 4   Column 12   Coefficient -0.03414154
         when "000000111100" => A <= "001101100011111111"; -- Line 4   Column 13   Coefficient 0.21191025
         when "000000111101" => A <= "000100010011001101"; -- Line 4   Column 14   Coefficient 0.06718826
         when "000000111110" => A <= "000000010111101010"; -- Line 4   Column 15   Coefficient 0.00577545
         when "000000111111" => A <= "111111111001000110"; -- Line 4   Column 16   Coefficient -0.00168610
         when "000001000000" => A <= "000000000000000110"; -- Line 5   Column 1   Coefficient 0.00002289
         when "000001000001" => A <= "000000000000000000"; -- Line 5   Column 2   Coefficient 0.00000000
         when "000001000010" => A <= "000000000000000000"; -- Line 5   Column 3   Coefficient 0.00000000
         when "000001000011" => A <= "000000000000000000"; -- Line 5   Column 4   Coefficient 0.00000000
         when "000001000100" => A <= "000000000000000000"; -- Line 5   Column 5   Coefficient 0.00000000
         when "000001000101" => A <= "000000000000000000"; -- Line 5   Column 6   Coefficient 0.00000000
         when "000001000110" => A <= "000000000000000000"; -- Line 5   Column 7   Coefficient 0.00000000
         when "000001000111" => A <= "000000000000000000"; -- Line 5   Column 8   Coefficient 0.00000000
         when "000001001000" => A <= "000000000000000000"; -- Line 5   Column 9   Coefficient 0.00000000
         when "000001001001" => A <= "000000000000000000"; -- Line 5   Column 10   Coefficient 0.00000000
         when "000001001010" => A <= "111111111111010011"; -- Line 5   Column 11   Coefficient -0.00017166
         when "000001001011" => A <= "111110000101010011"; -- Line 5   Column 12   Coefficient -0.02995682
         when "000001001100" => A <= "001100001011101000"; -- Line 5   Column 13   Coefficient 0.19033813
         when "000001001101" => A <= "000101100000010101"; -- Line 5   Column 14   Coefficient 0.08601761
         when "000001001110" => A <= "000000011000110111"; -- Line 5   Column 15   Coefficient 0.00606918
         when "000001001111" => A <= "111111110110011111"; -- Line 5   Column 16   Coefficient -0.00232315
         when "000001010000" => A <= "000000000000000100"; -- Line 6   Column 1   Coefficient 0.00001526
         when "000001010001" => A <= "000000000000000000"; -- Line 6   Column 2   Coefficient 0.00000000
         when "000001010010" => A <= "000000000000000000"; -- Line 6   Column 3   Coefficient 0.00000000
         when "000001010011" => A <= "000000000000000000"; -- Line 6   Column 4   Coefficient 0.00000000
         when "000001010100" => A <= "000000000000000000"; -- Line 6   Column 5   Coefficient 0.00000000
         when "000001010101" => A <= "000000000000000000"; -- Line 6   Column 6   Coefficient 0.00000000
         when "000001010110" => A <= "000000000000000000"; -- Line 6   Column 7   Coefficient 0.00000000
         when "000001010111" => A <= "000000000000000000"; -- Line 6   Column 8   Coefficient 0.00000000
         when "000001011000" => A <= "000000000000000000"; -- Line 6   Column 9   Coefficient 0.00000000
         when "000001011001" => A <= "000000000000000000"; -- Line 6   Column 10   Coefficient 0.00000000
         when "000001011010" => A <= "111111111110010010"; -- Line 6   Column 11   Coefficient -0.00041962
         when "000001011011" => A <= "111110010000110000"; -- Line 6   Column 12   Coefficient -0.02716064
         when "000001011100" => A <= "001010101100000111"; -- Line 6   Column 13   Coefficient 0.16701889
         when "000001011101" => A <= "000111000101010101"; -- Line 6   Column 14   Coefficient 0.11067581
         when "000001011110" => A <= "000000000100100100"; -- Line 6   Column 15   Coefficient 0.00111389
         when "000001011111" => A <= "111111111010111001"; -- Line 6   Column 16   Coefficient -0.00124741
         when "000001100000" => A <= "000000000000000011"; -- Line 7   Column 1   Coefficient 0.00001144
         when "000001100001" => A <= "000000000000000000"; -- Line 7   Column 2   Coefficient 0.00000000
         when "000001100010" => A <= "000000000000000000"; -- Line 7   Column 3   Coefficient 0.00000000
         when "000001100011" => A <= "000000000000000000"; -- Line 7   Column 4   Coefficient 0.00000000
         when "000001100100" => A <= "000000000000000000"; -- Line 7   Column 5   Coefficient 0.00000000
         when "000001100101" => A <= "000000000000000000"; -- Line 7   Column 6   Coefficient 0.00000000
         when "000001100110" => A <= "000000000000000000"; -- Line 7   Column 7   Coefficient 0.00000000
         when "000001100111" => A <= "000000000000000000"; -- Line 7   Column 8   Coefficient 0.00000000
         when "000001101000" => A <= "000000000000000000"; -- Line 7   Column 9   Coefficient 0.00000000
         when "000001101001" => A <= "000000000000000000"; -- Line 7   Column 10   Coefficient 0.00000000
         when "000001101010" => A <= "111111111110100110"; -- Line 7   Column 11   Coefficient -0.00034332
         when "000001101011" => A <= "111110011011111010"; -- Line 7   Column 12   Coefficient -0.02443695
         when "000001101100" => A <= "001001000110101001"; -- Line 7   Column 13   Coefficient 0.14224625
         when "000001101101" => A <= "001000110101000000"; -- Line 7   Column 14   Coefficient 0.13793945
         when "000001101110" => A <= "111111100111100010"; -- Line 7   Column 15   Coefficient -0.00597382
         when "000001101111" => A <= "000000000010010011"; -- Line 7   Column 16   Coefficient 0.00056076
         when "000001110000" => A <= "111111111111110100"; -- Line 8   Column 1   Coefficient -0.00004578
         when "000001110001" => A <= "000000000000000000"; -- Line 8   Column 2   Coefficient 0.00000000
         when "000001110010" => A <= "000000000000000000"; -- Line 8   Column 3   Coefficient 0.00000000
         when "000001110011" => A <= "000000000000000000"; -- Line 8   Column 4   Coefficient 0.00000000
         when "000001110100" => A <= "000000000000000000"; -- Line 8   Column 5   Coefficient 0.00000000
         when "000001110101" => A <= "000000000000000000"; -- Line 8   Column 6   Coefficient 0.00000000
         when "000001110110" => A <= "000000000000000000"; -- Line 8   Column 7   Coefficient 0.00000000
         when "000001110111" => A <= "000000000000000000"; -- Line 8   Column 8   Coefficient 0.00000000
         when "000001111000" => A <= "000000000000000000"; -- Line 8   Column 9   Coefficient 0.00000000
         when "000001111001" => A <= "000000000000000000"; -- Line 8   Column 10   Coefficient 0.00000000
         when "000001111010" => A <= "111111111111001011"; -- Line 8   Column 11   Coefficient -0.00020218
         when "000001111011" => A <= "111110100110010011"; -- Line 8   Column 12   Coefficient -0.02190018
         when "000001111100" => A <= "000111100110110001"; -- Line 8   Column 13   Coefficient 0.11883926
         when "000001111101" => A <= "001010011001111000"; -- Line 8   Column 14   Coefficient 0.16256714
         when "000001111110" => A <= "111111010000101110"; -- Line 8   Column 15   Coefficient -0.01154327
         when "000001111111" => A <= "000000001001011000"; -- Line 8   Column 16   Coefficient 0.00228882
         when "000010000000" => A <= "111111111111100110"; -- Line 9   Column 1   Coefficient -0.00009918
         when "000010000001" => A <= "000000000000000000"; -- Line 9   Column 2   Coefficient 0.00000000
         when "000010000010" => A <= "000000000000000000"; -- Line 9   Column 3   Coefficient 0.00000000
         when "000010000011" => A <= "000000000000000000"; -- Line 9   Column 4   Coefficient 0.00000000
         when "000010000100" => A <= "000000000000000000"; -- Line 9   Column 5   Coefficient 0.00000000
         when "000010000101" => A <= "000000000000000000"; -- Line 9   Column 6   Coefficient 0.00000000
         when "000010000110" => A <= "000000000000000000"; -- Line 9   Column 7   Coefficient 0.00000000
         when "000010000111" => A <= "000000000000000000"; -- Line 9   Column 8   Coefficient 0.00000000
         when "000010001000" => A <= "000000000000000000"; -- Line 9   Column 9   Coefficient 0.00000000
         when "000010001001" => A <= "000000000000000000"; -- Line 9   Column 10   Coefficient 0.00000000
         when "000010001010" => A <= "000000000000000011"; -- Line 9   Column 11   Coefficient 0.00001144
         when "000010001011" => A <= "111110110001100001"; -- Line 9   Column 12   Coefficient -0.01916122
         when "000010001100" => A <= "000110000101110011"; -- Line 9   Column 13   Coefficient 0.09516525
         when "000010001101" => A <= "001011111101111010"; -- Line 9   Column 14   Coefficient 0.18698883
         when "000010001110" => A <= "111110111010000001"; -- Line 9   Column 15   Coefficient -0.01708603
         when "000010001111" => A <= "000000010001001000"; -- Line 9   Column 16   Coefficient 0.00418091
         when "000010010000" => A <= "000000000000000111"; -- Line 10   Column 1   Coefficient 0.00002670
         when "000010010001" => A <= "000000000000000000"; -- Line 10   Column 2   Coefficient 0.00000000
         when "000010010010" => A <= "000000000000000000"; -- Line 10   Column 3   Coefficient 0.00000000
         when "000010010011" => A <= "000000000000000000"; -- Line 10   Column 4   Coefficient 0.00000000
         when "000010010100" => A <= "000000000000000000"; -- Line 10   Column 5   Coefficient 0.00000000
         when "000010010101" => A <= "000000000000000000"; -- Line 10   Column 6   Coefficient 0.00000000
         when "000010010110" => A <= "000000000000000000"; -- Line 10   Column 7   Coefficient 0.00000000
         when "000010010111" => A <= "000000000000000000"; -- Line 10   Column 8   Coefficient 0.00000000
         when "000010011000" => A <= "000000000000000000"; -- Line 10   Column 9   Coefficient 0.00000000
         when "000010011001" => A <= "000000000000000000"; -- Line 10   Column 10   Coefficient 0.00000000
         when "000010011010" => A <= "000000000000001001"; -- Line 10   Column 11   Coefficient 0.00003433
         when "000010011011" => A <= "111111000100111001"; -- Line 10   Column 12   Coefficient -0.01443100
         when "000010011100" => A <= "000100010010000101"; -- Line 10   Column 13   Coefficient 0.06691360
         when "000010011101" => A <= "001101110100101001"; -- Line 10   Column 14   Coefficient 0.21597672
         when "000010011110" => A <= "111110011010010101"; -- Line 10   Column 15   Coefficient -0.02482224
         when "000010011111" => A <= "000000011001110100"; -- Line 10   Column 16   Coefficient 0.00630188
         when "000010100000" => A <= "000000000000110011"; -- Line 11   Column 1   Coefficient 0.00019455
         when "000010100001" => A <= "000000000000000000"; -- Line 11   Column 2   Coefficient 0.00000000
         when "000010100010" => A <= "000000000000000000"; -- Line 11   Column 3   Coefficient 0.00000000
         when "000010100011" => A <= "000000000000000000"; -- Line 11   Column 4   Coefficient 0.00000000
         when "000010100100" => A <= "000000000000000000"; -- Line 11   Column 5   Coefficient 0.00000000
         when "000010100101" => A <= "000000000000000000"; -- Line 11   Column 6   Coefficient 0.00000000
         when "000010100110" => A <= "000000000000000000"; -- Line 11   Column 7   Coefficient 0.00000000
         when "000010100111" => A <= "000000000000000000"; -- Line 11   Column 8   Coefficient 0.00000000
         when "000010101000" => A <= "000000000000000000"; -- Line 11   Column 9   Coefficient 0.00000000
         when "000010101001" => A <= "000000000000000000"; -- Line 11   Column 10   Coefficient 0.00000000
         when "000010101010" => A <= "000000000000000000"; -- Line 11   Column 11   Coefficient 0.00000000
         when "000010101011" => A <= "111111011001111001"; -- Line 11   Column 12   Coefficient -0.00930405
         when "000010101100" => A <= "000010011110111100"; -- Line 11   Column 13   Coefficient 0.03880310
         when "000010101101" => A <= "001111100101110011"; -- Line 11   Column 14   Coefficient 0.24360275
         when "000010101110" => A <= "111101111110110001"; -- Line 11   Column 15   Coefficient -0.03155136
         when "000010101111" => A <= "000000100001110011"; -- Line 11   Column 16   Coefficient 0.00825119
         when "000010110000" => A <= "000000000001100101"; -- Line 12   Column 1   Coefficient 0.00038528
         when "000010110001" => A <= "000000000000000000"; -- Line 12   Column 2   Coefficient 0.00000000
         when "000010110010" => A <= "000000000000000000"; -- Line 12   Column 3   Coefficient 0.00000000
         when "000010110011" => A <= "000000000000000000"; -- Line 12   Column 4   Coefficient 0.00000000
         when "000010110100" => A <= "000000000000000000"; -- Line 12   Column 5   Coefficient 0.00000000
         when "000010110101" => A <= "000000000000000000"; -- Line 12   Column 6   Coefficient 0.00000000
         when "000010110110" => A <= "000000000000000000"; -- Line 12   Column 7   Coefficient 0.00000000
         when "000010110111" => A <= "000000000000000000"; -- Line 12   Column 8   Coefficient 0.00000000
         when "000010111000" => A <= "000000000000000000"; -- Line 12   Column 9   Coefficient 0.00000000
         when "000010111001" => A <= "000000000000000000"; -- Line 12   Column 10   Coefficient 0.00000000
         when "000010111010" => A <= "000000000000000000"; -- Line 12   Column 11   Coefficient 0.00000000
         when "000010111011" => A <= "111111110001010101"; -- Line 12   Column 12   Coefficient -0.00358200
         when "000010111100" => A <= "000000100101011001"; -- Line 12   Column 13   Coefficient 0.00912857
         when "000010111101" => A <= "010001011110001011"; -- Line 12   Column 14   Coefficient 0.27299118
         when "000010111110" => A <= "111101011101101101"; -- Line 12   Column 15   Coefficient -0.03962326
         when "000010111111" => A <= "000000101011110101"; -- Line 12   Column 16   Coefficient 0.01070023
         when "000011000000" => A <= "000000000010010101"; -- Line 13   Column 1   Coefficient 0.00056839
         when "000011000001" => A <= "000000000000000000"; -- Line 13   Column 2   Coefficient 0.00000000
         when "000011000010" => A <= "000000000000000000"; -- Line 13   Column 3   Coefficient 0.00000000
         when "000011000011" => A <= "000000000000000000"; -- Line 13   Column 4   Coefficient 0.00000000
         when "000011000100" => A <= "000000000000000000"; -- Line 13   Column 5   Coefficient 0.00000000
         when "000011000101" => A <= "000000000000000000"; -- Line 13   Column 6   Coefficient 0.00000000
         when "000011000110" => A <= "000000000000000000"; -- Line 13   Column 7   Coefficient 0.00000000
         when "000011000111" => A <= "000000000000000000"; -- Line 13   Column 8   Coefficient 0.00000000
         when "000011001000" => A <= "000000000000000000"; -- Line 13   Column 9   Coefficient 0.00000000
         when "000011001001" => A <= "000000000000000000"; -- Line 13   Column 10   Coefficient 0.00000000
         when "000011001010" => A <= "000000000000000000"; -- Line 13   Column 11   Coefficient 0.00000000
         when "000011001011" => A <= "000000000111011010"; -- Line 13   Column 12   Coefficient 0.00180817
         when "000011001100" => A <= "111110110101100100"; -- Line 13   Column 13   Coefficient -0.01817322
         when "000011001101" => A <= "010011000101100111"; -- Line 13   Column 14   Coefficient 0.29824448
         when "000011001110" => A <= "111101000110110001"; -- Line 13   Column 15   Coefficient -0.04522324
         when "000011001111" => A <= "000000110100010110"; -- Line 13   Column 16   Coefficient 0.01277924
         when "000011010000" => A <= "000000000001111110"; -- Line 14   Column 1   Coefficient 0.00048065
         when "000011010001" => A <= "000000000000000000"; -- Line 14   Column 2   Coefficient 0.00000000
         when "000011010010" => A <= "000000000000000000"; -- Line 14   Column 3   Coefficient 0.00000000
         when "000011010011" => A <= "000000000000000000"; -- Line 14   Column 4   Coefficient 0.00000000
         when "000011010100" => A <= "000000000000000000"; -- Line 14   Column 5   Coefficient 0.00000000
         when "000011010101" => A <= "000000000000000000"; -- Line 14   Column 6   Coefficient 0.00000000
         when "000011010110" => A <= "000000000000000000"; -- Line 14   Column 7   Coefficient 0.00000000
         when "000011010111" => A <= "000000000000000000"; -- Line 14   Column 8   Coefficient 0.00000000
         when "000011011000" => A <= "000000000000000000"; -- Line 14   Column 9   Coefficient 0.00000000
         when "000011011001" => A <= "000000000000000000"; -- Line 14   Column 10   Coefficient 0.00000000
         when "000011011010" => A <= "000000000000000000"; -- Line 14   Column 11   Coefficient 0.00000000
         when "000011011011" => A <= "000000001111000010"; -- Line 14   Column 12   Coefficient 0.00366974
         when "000011011100" => A <= "111110000010011110"; -- Line 14   Column 13   Coefficient -0.03064728
         when "000011011101" => A <= "010011010010100110"; -- Line 14   Column 14   Coefficient 0.30141449
         when "000011011110" => A <= "111101100111001110"; -- Line 14   Column 15   Coefficient -0.03730011
         when "000011011111" => A <= "000000110010101110"; -- Line 14   Column 16   Coefficient 0.01238251
         when "000011100000" => A <= "000000000001000010"; -- Line 15   Column 1   Coefficient 0.00025177
         when "000011100001" => A <= "000000000000000000"; -- Line 15   Column 2   Coefficient 0.00000000
         when "000011100010" => A <= "000000000000000000"; -- Line 15   Column 3   Coefficient 0.00000000
         when "000011100011" => A <= "000000000000000000"; -- Line 15   Column 4   Coefficient 0.00000000
         when "000011100100" => A <= "000000000000000000"; -- Line 15   Column 5   Coefficient 0.00000000
         when "000011100101" => A <= "000000000000000000"; -- Line 15   Column 6   Coefficient 0.00000000
         when "000011100110" => A <= "000000000000000000"; -- Line 15   Column 7   Coefficient 0.00000000
         when "000011100111" => A <= "000000000000000000"; -- Line 15   Column 8   Coefficient 0.00000000
         when "000011101000" => A <= "000000000000000000"; -- Line 15   Column 9   Coefficient 0.00000000
         when "000011101001" => A <= "000000000000000000"; -- Line 15   Column 10   Coefficient 0.00000000
         when "000011101010" => A <= "000000000000000000"; -- Line 15   Column 11   Coefficient 0.00000000
         when "000011101011" => A <= "000000010000011000"; -- Line 15   Column 12   Coefficient 0.00399780
         when "000011101100" => A <= "111101101011101110"; -- Line 15   Column 13   Coefficient -0.03620148
         when "000011101101" => A <= "010010110100110100"; -- Line 15   Column 14   Coefficient 0.29414368
         when "000011101110" => A <= "111110100000101100"; -- Line 15   Column 15   Coefficient -0.02326965
         when "000011101111" => A <= "000000101101010111"; -- Line 15   Column 16   Coefficient 0.01107407
         when "000011110000" => A <= "000000000001001000"; -- Line 16   Column 1   Coefficient 0.00027466
         when "000011110001" => A <= "000000000000000000"; -- Line 16   Column 2   Coefficient 0.00000000
         when "000011110010" => A <= "000000000000000000"; -- Line 16   Column 3   Coefficient 0.00000000
         when "000011110011" => A <= "000000000000000000"; -- Line 16   Column 4   Coefficient 0.00000000
         when "000011110100" => A <= "000000000000000000"; -- Line 16   Column 5   Coefficient 0.00000000
         when "000011110101" => A <= "000000000000000000"; -- Line 16   Column 6   Coefficient 0.00000000
         when "000011110110" => A <= "000000000000000000"; -- Line 16   Column 7   Coefficient 0.00000000
         when "000011110111" => A <= "000000000000000000"; -- Line 16   Column 8   Coefficient 0.00000000
         when "000011111000" => A <= "000000000000000000"; -- Line 16   Column 9   Coefficient 0.00000000
         when "000011111001" => A <= "000000000000000000"; -- Line 16   Column 10   Coefficient 0.00000000
         when "000011111010" => A <= "000000000000000000"; -- Line 16   Column 11   Coefficient 0.00000000
         when "000011111011" => A <= "000000001111111100"; -- Line 16   Column 12   Coefficient 0.00389099
         when "000011111100" => A <= "111101100000101101"; -- Line 16   Column 13   Coefficient -0.03889084
         when "000011111101" => A <= "010010000001100011"; -- Line 16   Column 14   Coefficient 0.28162766
         when "000011111110" => A <= "111111101010001000"; -- Line 16   Column 15   Coefficient -0.00534058
         when "000011111111" => A <= "000000100010100100"; -- Line 16   Column 16   Coefficient 0.00843811
         when "000100000000" => A <= "000000000001001011"; -- Line 17   Column 1   Coefficient 0.00028610
         when "000100000001" => A <= "000000000000000000"; -- Line 17   Column 2   Coefficient 0.00000000
         when "000100000010" => A <= "000000000000000000"; -- Line 17   Column 3   Coefficient 0.00000000
         when "000100000011" => A <= "000000000000000000"; -- Line 17   Column 4   Coefficient 0.00000000
         when "000100000100" => A <= "000000000000000000"; -- Line 17   Column 5   Coefficient 0.00000000
         when "000100000101" => A <= "000000000000000000"; -- Line 17   Column 6   Coefficient 0.00000000
         when "000100000110" => A <= "000000000000000000"; -- Line 17   Column 7   Coefficient 0.00000000
         when "000100000111" => A <= "000000000000000000"; -- Line 17   Column 8   Coefficient 0.00000000
         when "000100001000" => A <= "000000000000000000"; -- Line 17   Column 9   Coefficient 0.00000000
         when "000100001001" => A <= "000000000000000000"; -- Line 17   Column 10   Coefficient 0.00000000
         when "000100001010" => A <= "000000000000000000"; -- Line 17   Column 11   Coefficient 0.00000000
         when "000100001011" => A <= "000000001101001100"; -- Line 17   Column 12   Coefficient 0.00321960
         when "000100001100" => A <= "111101100010001110"; -- Line 17   Column 13   Coefficient -0.03852081
         when "000100001101" => A <= "010000111010100101"; -- Line 17   Column 14   Coefficient 0.26430130
         when "000100001110" => A <= "000000111110100110"; -- Line 17   Column 15   Coefficient 0.01528168
         when "000100001111" => A <= "000000010110010000"; -- Line 17   Column 16   Coefficient 0.00543213
         when "000100010000" => A <= "111111111110110111"; -- Line 18   Column 1   Coefficient -0.00027847
         when "000100010001" => A <= "000000000000000000"; -- Line 18   Column 2   Coefficient 0.00000000
         when "000100010010" => A <= "000000000000000000"; -- Line 18   Column 3   Coefficient 0.00000000
         when "000100010011" => A <= "000000000000000000"; -- Line 18   Column 4   Coefficient 0.00000000
         when "000100010100" => A <= "000000000000000000"; -- Line 18   Column 5   Coefficient 0.00000000
         when "000100010101" => A <= "000000000000000000"; -- Line 18   Column 6   Coefficient 0.00000000
         when "000100010110" => A <= "000000000000000000"; -- Line 18   Column 7   Coefficient 0.00000000
         when "000100010111" => A <= "000000000000000000"; -- Line 18   Column 8   Coefficient 0.00000000
         when "000100011000" => A <= "000000000000000000"; -- Line 18   Column 9   Coefficient 0.00000000
         when "000100011001" => A <= "000000000000000000"; -- Line 18   Column 10   Coefficient 0.00000000
         when "000100011010" => A <= "000000000000000000"; -- Line 18   Column 11   Coefficient 0.00000000
         when "000100011011" => A <= "000000001010110110"; -- Line 18   Column 12   Coefficient 0.00264740
         when "000100011100" => A <= "111101100010101111"; -- Line 18   Column 13   Coefficient -0.03839493
         when "000100011101" => A <= "001111111010100001"; -- Line 18   Column 14   Coefficient 0.24866104
         when "000100011110" => A <= "000010000100001011"; -- Line 18   Column 15   Coefficient 0.03226852
         when "000100011111" => A <= "000000010100110111"; -- Line 18   Column 16   Coefficient 0.00509262
         when "000100100000" => A <= "111111111100011110"; -- Line 19   Column 1   Coefficient -0.00086212
         when "000100100001" => A <= "111111111111111111"; -- Line 19   Column 2   Coefficient -0.00000381
         when "000100100010" => A <= "000000000000000000"; -- Line 19   Column 3   Coefficient 0.00000000
         when "000100100011" => A <= "000000000000000000"; -- Line 19   Column 4   Coefficient 0.00000000
         when "000100100100" => A <= "000000000000000000"; -- Line 19   Column 5   Coefficient 0.00000000
         when "000100100101" => A <= "000000000000000000"; -- Line 19   Column 6   Coefficient 0.00000000
         when "000100100110" => A <= "000000000000000000"; -- Line 19   Column 7   Coefficient 0.00000000
         when "000100100111" => A <= "000000000000000000"; -- Line 19   Column 8   Coefficient 0.00000000
         when "000100101000" => A <= "000000000000000000"; -- Line 19   Column 9   Coefficient 0.00000000
         when "000100101001" => A <= "000000000000000000"; -- Line 19   Column 10   Coefficient 0.00000000
         when "000100101010" => A <= "000000000000000000"; -- Line 19   Column 11   Coefficient 0.00000000
         when "000100101011" => A <= "000000001000010011"; -- Line 19   Column 12   Coefficient 0.00202560
         when "000100101100" => A <= "111101100110110000"; -- Line 19   Column 13   Coefficient -0.03741455
         when "000100101101" => A <= "001110110101010100"; -- Line 19   Column 14   Coefficient 0.23176575
         when "000100101110" => A <= "000011001010010011"; -- Line 19   Column 15   Coefficient 0.04938889
         when "000100101111" => A <= "000000010100111001"; -- Line 19   Column 16   Coefficient 0.00510025
         when "000100110000" => A <= "111111111001000110"; -- Line 20   Column 1   Coefficient -0.00168610
         when "000100110001" => A <= "000000000000000011"; -- Line 20   Column 2   Coefficient 0.00001144
         when "000100110010" => A <= "000000000000000000"; -- Line 20   Column 3   Coefficient 0.00000000
         when "000100110011" => A <= "000000000000000000"; -- Line 20   Column 4   Coefficient 0.00000000
         when "000100110100" => A <= "000000000000000000"; -- Line 20   Column 5   Coefficient 0.00000000
         when "000100110101" => A <= "000000000000000000"; -- Line 20   Column 6   Coefficient 0.00000000
         when "000100110110" => A <= "000000000000000000"; -- Line 20   Column 7   Coefficient 0.00000000
         when "000100110111" => A <= "000000000000000000"; -- Line 20   Column 8   Coefficient 0.00000000
         when "000100111000" => A <= "000000000000000000"; -- Line 20   Column 9   Coefficient 0.00000000
         when "000100111001" => A <= "000000000000000000"; -- Line 20   Column 10   Coefficient 0.00000000
         when "000100111010" => A <= "000000000000000000"; -- Line 20   Column 11   Coefficient 0.00000000
         when "000100111011" => A <= "000000000011111000"; -- Line 20   Column 12   Coefficient 0.00094604
         when "000100111100" => A <= "111101110100001010"; -- Line 20   Column 13   Coefficient -0.03414154
         when "000100111101" => A <= "001101100011111111"; -- Line 20   Column 14   Coefficient 0.21191025
         when "000100111110" => A <= "000100010011001101"; -- Line 20   Column 15   Coefficient 0.06718826
         when "000100111111" => A <= "000000010111101010"; -- Line 20   Column 16   Coefficient 0.00577545
         when "000101000000" => A <= "111111110110011111"; -- Line 21   Column 1   Coefficient -0.00232315
         when "000101000001" => A <= "000000000000000110"; -- Line 21   Column 2   Coefficient 0.00002289
         when "000101000010" => A <= "000000000000000000"; -- Line 21   Column 3   Coefficient 0.00000000
         when "000101000011" => A <= "000000000000000000"; -- Line 21   Column 4   Coefficient 0.00000000
         when "000101000100" => A <= "000000000000000000"; -- Line 21   Column 5   Coefficient 0.00000000
         when "000101000101" => A <= "000000000000000000"; -- Line 21   Column 6   Coefficient 0.00000000
         when "000101000110" => A <= "000000000000000000"; -- Line 21   Column 7   Coefficient 0.00000000
         when "000101000111" => A <= "000000000000000000"; -- Line 21   Column 8   Coefficient 0.00000000
         when "000101001000" => A <= "000000000000000000"; -- Line 21   Column 9   Coefficient 0.00000000
         when "000101001001" => A <= "000000000000000000"; -- Line 21   Column 10   Coefficient 0.00000000
         when "000101001010" => A <= "000000000000000000"; -- Line 21   Column 11   Coefficient 0.00000000
         when "000101001011" => A <= "111111111111010011"; -- Line 21   Column 12   Coefficient -0.00017166
         when "000101001100" => A <= "111110000101010011"; -- Line 21   Column 13   Coefficient -0.02995682
         when "000101001101" => A <= "001100001011101000"; -- Line 21   Column 14   Coefficient 0.19033813
         when "000101001110" => A <= "000101100000010101"; -- Line 21   Column 15   Coefficient 0.08601761
         when "000101001111" => A <= "000000011000110111"; -- Line 21   Column 16   Coefficient 0.00606918
         when "000101010000" => A <= "111111111010111001"; -- Line 22   Column 1   Coefficient -0.00124741
         when "000101010001" => A <= "000000000000000100"; -- Line 22   Column 2   Coefficient 0.00001526
         when "000101010010" => A <= "000000000000000000"; -- Line 22   Column 3   Coefficient 0.00000000
         when "000101010011" => A <= "000000000000000000"; -- Line 22   Column 4   Coefficient 0.00000000
         when "000101010100" => A <= "000000000000000000"; -- Line 22   Column 5   Coefficient 0.00000000
         when "000101010101" => A <= "000000000000000000"; -- Line 22   Column 6   Coefficient 0.00000000
         when "000101010110" => A <= "000000000000000000"; -- Line 22   Column 7   Coefficient 0.00000000
         when "000101010111" => A <= "000000000000000000"; -- Line 22   Column 8   Coefficient 0.00000000
         when "000101011000" => A <= "000000000000000000"; -- Line 22   Column 9   Coefficient 0.00000000
         when "000101011001" => A <= "000000000000000000"; -- Line 22   Column 10   Coefficient 0.00000000
         when "000101011010" => A <= "000000000000000000"; -- Line 22   Column 11   Coefficient 0.00000000
         when "000101011011" => A <= "111111111110010010"; -- Line 22   Column 12   Coefficient -0.00041962
         when "000101011100" => A <= "111110010000110000"; -- Line 22   Column 13   Coefficient -0.02716064
         when "000101011101" => A <= "001010101100000111"; -- Line 22   Column 14   Coefficient 0.16701889
         when "000101011110" => A <= "000111000101010101"; -- Line 22   Column 15   Coefficient 0.11067581
         when "000101011111" => A <= "000000000100100100"; -- Line 22   Column 16   Coefficient 0.00111389
         when "000101100000" => A <= "000000000010010011"; -- Line 23   Column 1   Coefficient 0.00056076
         when "000101100001" => A <= "000000000000000011"; -- Line 23   Column 2   Coefficient 0.00001144
         when "000101100010" => A <= "000000000000000000"; -- Line 23   Column 3   Coefficient 0.00000000
         when "000101100011" => A <= "000000000000000000"; -- Line 23   Column 4   Coefficient 0.00000000
         when "000101100100" => A <= "000000000000000000"; -- Line 23   Column 5   Coefficient 0.00000000
         when "000101100101" => A <= "000000000000000000"; -- Line 23   Column 6   Coefficient 0.00000000
         when "000101100110" => A <= "000000000000000000"; -- Line 23   Column 7   Coefficient 0.00000000
         when "000101100111" => A <= "000000000000000000"; -- Line 23   Column 8   Coefficient 0.00000000
         when "000101101000" => A <= "000000000000000000"; -- Line 23   Column 9   Coefficient 0.00000000
         when "000101101001" => A <= "000000000000000000"; -- Line 23   Column 10   Coefficient 0.00000000
         when "000101101010" => A <= "000000000000000000"; -- Line 23   Column 11   Coefficient 0.00000000
         when "000101101011" => A <= "111111111110100110"; -- Line 23   Column 12   Coefficient -0.00034332
         when "000101101100" => A <= "111110011011111010"; -- Line 23   Column 13   Coefficient -0.02443695
         when "000101101101" => A <= "001001000110101001"; -- Line 23   Column 14   Coefficient 0.14224625
         when "000101101110" => A <= "001000110101000000"; -- Line 23   Column 15   Coefficient 0.13793945
         when "000101101111" => A <= "111111100111100010"; -- Line 23   Column 16   Coefficient -0.00597382
         when "000101110000" => A <= "000000001001011000"; -- Line 24   Column 1   Coefficient 0.00228882
         when "000101110001" => A <= "111111111111110100"; -- Line 24   Column 2   Coefficient -0.00004578
         when "000101110010" => A <= "000000000000000000"; -- Line 24   Column 3   Coefficient 0.00000000
         when "000101110011" => A <= "000000000000000000"; -- Line 24   Column 4   Coefficient 0.00000000
         when "000101110100" => A <= "000000000000000000"; -- Line 24   Column 5   Coefficient 0.00000000
         when "000101110101" => A <= "000000000000000000"; -- Line 24   Column 6   Coefficient 0.00000000
         when "000101110110" => A <= "000000000000000000"; -- Line 24   Column 7   Coefficient 0.00000000
         when "000101110111" => A <= "000000000000000000"; -- Line 24   Column 8   Coefficient 0.00000000
         when "000101111000" => A <= "000000000000000000"; -- Line 24   Column 9   Coefficient 0.00000000
         when "000101111001" => A <= "000000000000000000"; -- Line 24   Column 10   Coefficient 0.00000000
         when "000101111010" => A <= "000000000000000000"; -- Line 24   Column 11   Coefficient 0.00000000
         when "000101111011" => A <= "111111111111001011"; -- Line 24   Column 12   Coefficient -0.00020218
         when "000101111100" => A <= "111110100110010011"; -- Line 24   Column 13   Coefficient -0.02190018
         when "000101111101" => A <= "000111100110110001"; -- Line 24   Column 14   Coefficient 0.11883926
         when "000101111110" => A <= "001010011001111000"; -- Line 24   Column 15   Coefficient 0.16256714
         when "000101111111" => A <= "111111010000101110"; -- Line 24   Column 16   Coefficient -0.01154327
         when "000110000000" => A <= "000000010001001000"; -- Line 25   Column 1   Coefficient 0.00418091
         when "000110000001" => A <= "111111111111100110"; -- Line 25   Column 2   Coefficient -0.00009918
         when "000110000010" => A <= "000000000000000000"; -- Line 25   Column 3   Coefficient 0.00000000
         when "000110000011" => A <= "000000000000000000"; -- Line 25   Column 4   Coefficient 0.00000000
         when "000110000100" => A <= "000000000000000000"; -- Line 25   Column 5   Coefficient 0.00000000
         when "000110000101" => A <= "000000000000000000"; -- Line 25   Column 6   Coefficient 0.00000000
         when "000110000110" => A <= "000000000000000000"; -- Line 25   Column 7   Coefficient 0.00000000
         when "000110000111" => A <= "000000000000000000"; -- Line 25   Column 8   Coefficient 0.00000000
         when "000110001000" => A <= "000000000000000000"; -- Line 25   Column 9   Coefficient 0.00000000
         when "000110001001" => A <= "000000000000000000"; -- Line 25   Column 10   Coefficient 0.00000000
         when "000110001010" => A <= "000000000000000000"; -- Line 25   Column 11   Coefficient 0.00000000
         when "000110001011" => A <= "000000000000000011"; -- Line 25   Column 12   Coefficient 0.00001144
         when "000110001100" => A <= "111110110001100001"; -- Line 25   Column 13   Coefficient -0.01916122
         when "000110001101" => A <= "000110000101110011"; -- Line 25   Column 14   Coefficient 0.09516525
         when "000110001110" => A <= "001011111101111010"; -- Line 25   Column 15   Coefficient 0.18698883
         when "000110001111" => A <= "111110111010000001"; -- Line 25   Column 16   Coefficient -0.01708603
         when "000110010000" => A <= "000000011001110100"; -- Line 26   Column 1   Coefficient 0.00630188
         when "000110010001" => A <= "000000000000000111"; -- Line 26   Column 2   Coefficient 0.00002670
         when "000110010010" => A <= "000000000000000000"; -- Line 26   Column 3   Coefficient 0.00000000
         when "000110010011" => A <= "000000000000000000"; -- Line 26   Column 4   Coefficient 0.00000000
         when "000110010100" => A <= "000000000000000000"; -- Line 26   Column 5   Coefficient 0.00000000
         when "000110010101" => A <= "000000000000000000"; -- Line 26   Column 6   Coefficient 0.00000000
         when "000110010110" => A <= "000000000000000000"; -- Line 26   Column 7   Coefficient 0.00000000
         when "000110010111" => A <= "000000000000000000"; -- Line 26   Column 8   Coefficient 0.00000000
         when "000110011000" => A <= "000000000000000000"; -- Line 26   Column 9   Coefficient 0.00000000
         when "000110011001" => A <= "000000000000000000"; -- Line 26   Column 10   Coefficient 0.00000000
         when "000110011010" => A <= "000000000000000000"; -- Line 26   Column 11   Coefficient 0.00000000
         when "000110011011" => A <= "000000000000001001"; -- Line 26   Column 12   Coefficient 0.00003433
         when "000110011100" => A <= "111111000100111001"; -- Line 26   Column 13   Coefficient -0.01443100
         when "000110011101" => A <= "000100010010000101"; -- Line 26   Column 14   Coefficient 0.06691360
         when "000110011110" => A <= "001101110100101001"; -- Line 26   Column 15   Coefficient 0.21597672
         when "000110011111" => A <= "111110011010010101"; -- Line 26   Column 16   Coefficient -0.02482224
         when "000110100000" => A <= "000000100001110011"; -- Line 27   Column 1   Coefficient 0.00825119
         when "000110100001" => A <= "000000000000110011"; -- Line 27   Column 2   Coefficient 0.00019455
         when "000110100010" => A <= "000000000000000000"; -- Line 27   Column 3   Coefficient 0.00000000
         when "000110100011" => A <= "000000000000000000"; -- Line 27   Column 4   Coefficient 0.00000000
         when "000110100100" => A <= "000000000000000000"; -- Line 27   Column 5   Coefficient 0.00000000
         when "000110100101" => A <= "000000000000000000"; -- Line 27   Column 6   Coefficient 0.00000000
         when "000110100110" => A <= "000000000000000000"; -- Line 27   Column 7   Coefficient 0.00000000
         when "000110100111" => A <= "000000000000000000"; -- Line 27   Column 8   Coefficient 0.00000000
         when "000110101000" => A <= "000000000000000000"; -- Line 27   Column 9   Coefficient 0.00000000
         when "000110101001" => A <= "000000000000000000"; -- Line 27   Column 10   Coefficient 0.00000000
         when "000110101010" => A <= "000000000000000000"; -- Line 27   Column 11   Coefficient 0.00000000
         when "000110101011" => A <= "000000000000000000"; -- Line 27   Column 12   Coefficient 0.00000000
         when "000110101100" => A <= "111111011001111001"; -- Line 27   Column 13   Coefficient -0.00930405
         when "000110101101" => A <= "000010011110111100"; -- Line 27   Column 14   Coefficient 0.03880310
         when "000110101110" => A <= "001111100101110011"; -- Line 27   Column 15   Coefficient 0.24360275
         when "000110101111" => A <= "111101111110110001"; -- Line 27   Column 16   Coefficient -0.03155136
         when "000110110000" => A <= "000000101011110101"; -- Line 28   Column 1   Coefficient 0.01070023
         when "000110110001" => A <= "000000000001100101"; -- Line 28   Column 2   Coefficient 0.00038528
         when "000110110010" => A <= "000000000000000000"; -- Line 28   Column 3   Coefficient 0.00000000
         when "000110110011" => A <= "000000000000000000"; -- Line 28   Column 4   Coefficient 0.00000000
         when "000110110100" => A <= "000000000000000000"; -- Line 28   Column 5   Coefficient 0.00000000
         when "000110110101" => A <= "000000000000000000"; -- Line 28   Column 6   Coefficient 0.00000000
         when "000110110110" => A <= "000000000000000000"; -- Line 28   Column 7   Coefficient 0.00000000
         when "000110110111" => A <= "000000000000000000"; -- Line 28   Column 8   Coefficient 0.00000000
         when "000110111000" => A <= "000000000000000000"; -- Line 28   Column 9   Coefficient 0.00000000
         when "000110111001" => A <= "000000000000000000"; -- Line 28   Column 10   Coefficient 0.00000000
         when "000110111010" => A <= "000000000000000000"; -- Line 28   Column 11   Coefficient 0.00000000
         when "000110111011" => A <= "000000000000000000"; -- Line 28   Column 12   Coefficient 0.00000000
         when "000110111100" => A <= "111111110001010101"; -- Line 28   Column 13   Coefficient -0.00358200
         when "000110111101" => A <= "000000100101011001"; -- Line 28   Column 14   Coefficient 0.00912857
         when "000110111110" => A <= "010001011110001011"; -- Line 28   Column 15   Coefficient 0.27299118
         when "000110111111" => A <= "111101011101101101"; -- Line 28   Column 16   Coefficient -0.03962326
         when "000111000000" => A <= "000000110100010110"; -- Line 29   Column 1   Coefficient 0.01277924
         when "000111000001" => A <= "000000000010010101"; -- Line 29   Column 2   Coefficient 0.00056839
         when "000111000010" => A <= "000000000000000000"; -- Line 29   Column 3   Coefficient 0.00000000
         when "000111000011" => A <= "000000000000000000"; -- Line 29   Column 4   Coefficient 0.00000000
         when "000111000100" => A <= "000000000000000000"; -- Line 29   Column 5   Coefficient 0.00000000
         when "000111000101" => A <= "000000000000000000"; -- Line 29   Column 6   Coefficient 0.00000000
         when "000111000110" => A <= "000000000000000000"; -- Line 29   Column 7   Coefficient 0.00000000
         when "000111000111" => A <= "000000000000000000"; -- Line 29   Column 8   Coefficient 0.00000000
         when "000111001000" => A <= "000000000000000000"; -- Line 29   Column 9   Coefficient 0.00000000
         when "000111001001" => A <= "000000000000000000"; -- Line 29   Column 10   Coefficient 0.00000000
         when "000111001010" => A <= "000000000000000000"; -- Line 29   Column 11   Coefficient 0.00000000
         when "000111001011" => A <= "000000000000000000"; -- Line 29   Column 12   Coefficient 0.00000000
         when "000111001100" => A <= "000000000111011010"; -- Line 29   Column 13   Coefficient 0.00180817
         when "000111001101" => A <= "111110110101100100"; -- Line 29   Column 14   Coefficient -0.01817322
         when "000111001110" => A <= "010011000101100111"; -- Line 29   Column 15   Coefficient 0.29824448
         when "000111001111" => A <= "111101000110110001"; -- Line 29   Column 16   Coefficient -0.04522324
         when "000111010000" => A <= "000000110010101110"; -- Line 30   Column 1   Coefficient 0.01238251
         when "000111010001" => A <= "000000000001111110"; -- Line 30   Column 2   Coefficient 0.00048065
         when "000111010010" => A <= "000000000000000000"; -- Line 30   Column 3   Coefficient 0.00000000
         when "000111010011" => A <= "000000000000000000"; -- Line 30   Column 4   Coefficient 0.00000000
         when "000111010100" => A <= "000000000000000000"; -- Line 30   Column 5   Coefficient 0.00000000
         when "000111010101" => A <= "000000000000000000"; -- Line 30   Column 6   Coefficient 0.00000000
         when "000111010110" => A <= "000000000000000000"; -- Line 30   Column 7   Coefficient 0.00000000
         when "000111010111" => A <= "000000000000000000"; -- Line 30   Column 8   Coefficient 0.00000000
         when "000111011000" => A <= "000000000000000000"; -- Line 30   Column 9   Coefficient 0.00000000
         when "000111011001" => A <= "000000000000000000"; -- Line 30   Column 10   Coefficient 0.00000000
         when "000111011010" => A <= "000000000000000000"; -- Line 30   Column 11   Coefficient 0.00000000
         when "000111011011" => A <= "000000000000000000"; -- Line 30   Column 12   Coefficient 0.00000000
         when "000111011100" => A <= "000000001111000010"; -- Line 30   Column 13   Coefficient 0.00366974
         when "000111011101" => A <= "111110000010011110"; -- Line 30   Column 14   Coefficient -0.03064728
         when "000111011110" => A <= "010011010010100110"; -- Line 30   Column 15   Coefficient 0.30141449
         when "000111011111" => A <= "111101100111001110"; -- Line 30   Column 16   Coefficient -0.03730011
         when "000111100000" => A <= "000000101101010111"; -- Line 31   Column 1   Coefficient 0.01107407
         when "000111100001" => A <= "000000000001000010"; -- Line 31   Column 2   Coefficient 0.00025177
         when "000111100010" => A <= "000000000000000000"; -- Line 31   Column 3   Coefficient 0.00000000
         when "000111100011" => A <= "000000000000000000"; -- Line 31   Column 4   Coefficient 0.00000000
         when "000111100100" => A <= "000000000000000000"; -- Line 31   Column 5   Coefficient 0.00000000
         when "000111100101" => A <= "000000000000000000"; -- Line 31   Column 6   Coefficient 0.00000000
         when "000111100110" => A <= "000000000000000000"; -- Line 31   Column 7   Coefficient 0.00000000
         when "000111100111" => A <= "000000000000000000"; -- Line 31   Column 8   Coefficient 0.00000000
         when "000111101000" => A <= "000000000000000000"; -- Line 31   Column 9   Coefficient 0.00000000
         when "000111101001" => A <= "000000000000000000"; -- Line 31   Column 10   Coefficient 0.00000000
         when "000111101010" => A <= "000000000000000000"; -- Line 31   Column 11   Coefficient 0.00000000
         when "000111101011" => A <= "000000000000000000"; -- Line 31   Column 12   Coefficient 0.00000000
         when "000111101100" => A <= "000000010000011000"; -- Line 31   Column 13   Coefficient 0.00399780
         when "000111101101" => A <= "111101101011101110"; -- Line 31   Column 14   Coefficient -0.03620148
         when "000111101110" => A <= "010010110100110100"; -- Line 31   Column 15   Coefficient 0.29414368
         when "000111101111" => A <= "111110100000101100"; -- Line 31   Column 16   Coefficient -0.02326965
         when "000111110000" => A <= "000000100010100100"; -- Line 32   Column 1   Coefficient 0.00843811
         when "000111110001" => A <= "000000000001001000"; -- Line 32   Column 2   Coefficient 0.00027466
         when "000111110010" => A <= "000000000000000000"; -- Line 32   Column 3   Coefficient 0.00000000
         when "000111110011" => A <= "000000000000000000"; -- Line 32   Column 4   Coefficient 0.00000000
         when "000111110100" => A <= "000000000000000000"; -- Line 32   Column 5   Coefficient 0.00000000
         when "000111110101" => A <= "000000000000000000"; -- Line 32   Column 6   Coefficient 0.00000000
         when "000111110110" => A <= "000000000000000000"; -- Line 32   Column 7   Coefficient 0.00000000
         when "000111110111" => A <= "000000000000000000"; -- Line 32   Column 8   Coefficient 0.00000000
         when "000111111000" => A <= "000000000000000000"; -- Line 32   Column 9   Coefficient 0.00000000
         when "000111111001" => A <= "000000000000000000"; -- Line 32   Column 10   Coefficient 0.00000000
         when "000111111010" => A <= "000000000000000000"; -- Line 32   Column 11   Coefficient 0.00000000
         when "000111111011" => A <= "000000000000000000"; -- Line 32   Column 12   Coefficient 0.00000000
         when "000111111100" => A <= "000000001111111100"; -- Line 32   Column 13   Coefficient 0.00389099
         when "000111111101" => A <= "111101100000101101"; -- Line 32   Column 14   Coefficient -0.03889084
         when "000111111110" => A <= "010010000001100011"; -- Line 32   Column 15   Coefficient 0.28162766
         when "000111111111" => A <= "111111101010001000"; -- Line 32   Column 16   Coefficient -0.00534058
         when "001000000000" => A <= "000000010110010000"; -- Line 33   Column 1   Coefficient 0.00543213
         when "001000000001" => A <= "000000000001001011"; -- Line 33   Column 2   Coefficient 0.00028610
         when "001000000010" => A <= "000000000000000000"; -- Line 33   Column 3   Coefficient 0.00000000
         when "001000000011" => A <= "000000000000000000"; -- Line 33   Column 4   Coefficient 0.00000000
         when "001000000100" => A <= "000000000000000000"; -- Line 33   Column 5   Coefficient 0.00000000
         when "001000000101" => A <= "000000000000000000"; -- Line 33   Column 6   Coefficient 0.00000000
         when "001000000110" => A <= "000000000000000000"; -- Line 33   Column 7   Coefficient 0.00000000
         when "001000000111" => A <= "000000000000000000"; -- Line 33   Column 8   Coefficient 0.00000000
         when "001000001000" => A <= "000000000000000000"; -- Line 33   Column 9   Coefficient 0.00000000
         when "001000001001" => A <= "000000000000000000"; -- Line 33   Column 10   Coefficient 0.00000000
         when "001000001010" => A <= "000000000000000000"; -- Line 33   Column 11   Coefficient 0.00000000
         when "001000001011" => A <= "000000000000000000"; -- Line 33   Column 12   Coefficient 0.00000000
         when "001000001100" => A <= "000000001101001100"; -- Line 33   Column 13   Coefficient 0.00321960
         when "001000001101" => A <= "111101100010001110"; -- Line 33   Column 14   Coefficient -0.03852081
         when "001000001110" => A <= "010000111010100101"; -- Line 33   Column 15   Coefficient 0.26430130
         when "001000001111" => A <= "000000111110100110"; -- Line 33   Column 16   Coefficient 0.01528168
         when "001000010000" => A <= "000000010100110111"; -- Line 34   Column 1   Coefficient 0.00509262
         when "001000010001" => A <= "111111111110110111"; -- Line 34   Column 2   Coefficient -0.00027847
         when "001000010010" => A <= "000000000000000000"; -- Line 34   Column 3   Coefficient 0.00000000
         when "001000010011" => A <= "000000000000000000"; -- Line 34   Column 4   Coefficient 0.00000000
         when "001000010100" => A <= "000000000000000000"; -- Line 34   Column 5   Coefficient 0.00000000
         when "001000010101" => A <= "000000000000000000"; -- Line 34   Column 6   Coefficient 0.00000000
         when "001000010110" => A <= "000000000000000000"; -- Line 34   Column 7   Coefficient 0.00000000
         when "001000010111" => A <= "000000000000000000"; -- Line 34   Column 8   Coefficient 0.00000000
         when "001000011000" => A <= "000000000000000000"; -- Line 34   Column 9   Coefficient 0.00000000
         when "001000011001" => A <= "000000000000000000"; -- Line 34   Column 10   Coefficient 0.00000000
         when "001000011010" => A <= "000000000000000000"; -- Line 34   Column 11   Coefficient 0.00000000
         when "001000011011" => A <= "000000000000000000"; -- Line 34   Column 12   Coefficient 0.00000000
         when "001000011100" => A <= "000000001010110110"; -- Line 34   Column 13   Coefficient 0.00264740
         when "001000011101" => A <= "111101100010101111"; -- Line 34   Column 14   Coefficient -0.03839493
         when "001000011110" => A <= "001111111010100001"; -- Line 34   Column 15   Coefficient 0.24866104
         when "001000011111" => A <= "000010000100001011"; -- Line 34   Column 16   Coefficient 0.03226852
         when "001000100000" => A <= "000000010100111001"; -- Line 35   Column 1   Coefficient 0.00510025
         when "001000100001" => A <= "111111111100011110"; -- Line 35   Column 2   Coefficient -0.00086212
         when "001000100010" => A <= "111111111111111111"; -- Line 35   Column 3   Coefficient -0.00000381
         when "001000100011" => A <= "000000000000000000"; -- Line 35   Column 4   Coefficient 0.00000000
         when "001000100100" => A <= "000000000000000000"; -- Line 35   Column 5   Coefficient 0.00000000
         when "001000100101" => A <= "000000000000000000"; -- Line 35   Column 6   Coefficient 0.00000000
         when "001000100110" => A <= "000000000000000000"; -- Line 35   Column 7   Coefficient 0.00000000
         when "001000100111" => A <= "000000000000000000"; -- Line 35   Column 8   Coefficient 0.00000000
         when "001000101000" => A <= "000000000000000000"; -- Line 35   Column 9   Coefficient 0.00000000
         when "001000101001" => A <= "000000000000000000"; -- Line 35   Column 10   Coefficient 0.00000000
         when "001000101010" => A <= "000000000000000000"; -- Line 35   Column 11   Coefficient 0.00000000
         when "001000101011" => A <= "000000000000000000"; -- Line 35   Column 12   Coefficient 0.00000000
         when "001000101100" => A <= "000000001000010011"; -- Line 35   Column 13   Coefficient 0.00202560
         when "001000101101" => A <= "111101100110110000"; -- Line 35   Column 14   Coefficient -0.03741455
         when "001000101110" => A <= "001110110101010100"; -- Line 35   Column 15   Coefficient 0.23176575
         when "001000101111" => A <= "000011001010010011"; -- Line 35   Column 16   Coefficient 0.04938889
         when "001000110000" => A <= "000000010111101010"; -- Line 36   Column 1   Coefficient 0.00577545
         when "001000110001" => A <= "111111111001000110"; -- Line 36   Column 2   Coefficient -0.00168610
         when "001000110010" => A <= "000000000000000011"; -- Line 36   Column 3   Coefficient 0.00001144
         when "001000110011" => A <= "000000000000000000"; -- Line 36   Column 4   Coefficient 0.00000000
         when "001000110100" => A <= "000000000000000000"; -- Line 36   Column 5   Coefficient 0.00000000
         when "001000110101" => A <= "000000000000000000"; -- Line 36   Column 6   Coefficient 0.00000000
         when "001000110110" => A <= "000000000000000000"; -- Line 36   Column 7   Coefficient 0.00000000
         when "001000110111" => A <= "000000000000000000"; -- Line 36   Column 8   Coefficient 0.00000000
         when "001000111000" => A <= "000000000000000000"; -- Line 36   Column 9   Coefficient 0.00000000
         when "001000111001" => A <= "000000000000000000"; -- Line 36   Column 10   Coefficient 0.00000000
         when "001000111010" => A <= "000000000000000000"; -- Line 36   Column 11   Coefficient 0.00000000
         when "001000111011" => A <= "000000000000000000"; -- Line 36   Column 12   Coefficient 0.00000000
         when "001000111100" => A <= "000000000011111000"; -- Line 36   Column 13   Coefficient 0.00094604
         when "001000111101" => A <= "111101110100001010"; -- Line 36   Column 14   Coefficient -0.03414154
         when "001000111110" => A <= "001101100011111111"; -- Line 36   Column 15   Coefficient 0.21191025
         when "001000111111" => A <= "000100010011001101"; -- Line 36   Column 16   Coefficient 0.06718826
         when "001001000000" => A <= "000000011000110111"; -- Line 37   Column 1   Coefficient 0.00606918
         when "001001000001" => A <= "111111110110011111"; -- Line 37   Column 2   Coefficient -0.00232315
         when "001001000010" => A <= "000000000000000110"; -- Line 37   Column 3   Coefficient 0.00002289
         when "001001000011" => A <= "000000000000000000"; -- Line 37   Column 4   Coefficient 0.00000000
         when "001001000100" => A <= "000000000000000000"; -- Line 37   Column 5   Coefficient 0.00000000
         when "001001000101" => A <= "000000000000000000"; -- Line 37   Column 6   Coefficient 0.00000000
         when "001001000110" => A <= "000000000000000000"; -- Line 37   Column 7   Coefficient 0.00000000
         when "001001000111" => A <= "000000000000000000"; -- Line 37   Column 8   Coefficient 0.00000000
         when "001001001000" => A <= "000000000000000000"; -- Line 37   Column 9   Coefficient 0.00000000
         when "001001001001" => A <= "000000000000000000"; -- Line 37   Column 10   Coefficient 0.00000000
         when "001001001010" => A <= "000000000000000000"; -- Line 37   Column 11   Coefficient 0.00000000
         when "001001001011" => A <= "000000000000000000"; -- Line 37   Column 12   Coefficient 0.00000000
         when "001001001100" => A <= "111111111111010011"; -- Line 37   Column 13   Coefficient -0.00017166
         when "001001001101" => A <= "111110000101010011"; -- Line 37   Column 14   Coefficient -0.02995682
         when "001001001110" => A <= "001100001011101000"; -- Line 37   Column 15   Coefficient 0.19033813
         when "001001001111" => A <= "000101100000010101"; -- Line 37   Column 16   Coefficient 0.08601761
         when "001001010000" => A <= "000000000100100100"; -- Line 38   Column 1   Coefficient 0.00111389
         when "001001010001" => A <= "111111111010111001"; -- Line 38   Column 2   Coefficient -0.00124741
         when "001001010010" => A <= "000000000000000100"; -- Line 38   Column 3   Coefficient 0.00001526
         when "001001010011" => A <= "000000000000000000"; -- Line 38   Column 4   Coefficient 0.00000000
         when "001001010100" => A <= "000000000000000000"; -- Line 38   Column 5   Coefficient 0.00000000
         when "001001010101" => A <= "000000000000000000"; -- Line 38   Column 6   Coefficient 0.00000000
         when "001001010110" => A <= "000000000000000000"; -- Line 38   Column 7   Coefficient 0.00000000
         when "001001010111" => A <= "000000000000000000"; -- Line 38   Column 8   Coefficient 0.00000000
         when "001001011000" => A <= "000000000000000000"; -- Line 38   Column 9   Coefficient 0.00000000
         when "001001011001" => A <= "000000000000000000"; -- Line 38   Column 10   Coefficient 0.00000000
         when "001001011010" => A <= "000000000000000000"; -- Line 38   Column 11   Coefficient 0.00000000
         when "001001011011" => A <= "000000000000000000"; -- Line 38   Column 12   Coefficient 0.00000000
         when "001001011100" => A <= "111111111110010010"; -- Line 38   Column 13   Coefficient -0.00041962
         when "001001011101" => A <= "111110010000110000"; -- Line 38   Column 14   Coefficient -0.02716064
         when "001001011110" => A <= "001010101100000111"; -- Line 38   Column 15   Coefficient 0.16701889
         when "001001011111" => A <= "000111000101010101"; -- Line 38   Column 16   Coefficient 0.11067581
         when "001001100000" => A <= "111111100111100010"; -- Line 39   Column 1   Coefficient -0.00597382
         when "001001100001" => A <= "000000000010010011"; -- Line 39   Column 2   Coefficient 0.00056076
         when "001001100010" => A <= "000000000000000011"; -- Line 39   Column 3   Coefficient 0.00001144
         when "001001100011" => A <= "000000000000000000"; -- Line 39   Column 4   Coefficient 0.00000000
         when "001001100100" => A <= "000000000000000000"; -- Line 39   Column 5   Coefficient 0.00000000
         when "001001100101" => A <= "000000000000000000"; -- Line 39   Column 6   Coefficient 0.00000000
         when "001001100110" => A <= "000000000000000000"; -- Line 39   Column 7   Coefficient 0.00000000
         when "001001100111" => A <= "000000000000000000"; -- Line 39   Column 8   Coefficient 0.00000000
         when "001001101000" => A <= "000000000000000000"; -- Line 39   Column 9   Coefficient 0.00000000
         when "001001101001" => A <= "000000000000000000"; -- Line 39   Column 10   Coefficient 0.00000000
         when "001001101010" => A <= "000000000000000000"; -- Line 39   Column 11   Coefficient 0.00000000
         when "001001101011" => A <= "000000000000000000"; -- Line 39   Column 12   Coefficient 0.00000000
         when "001001101100" => A <= "111111111110100110"; -- Line 39   Column 13   Coefficient -0.00034332
         when "001001101101" => A <= "111110011011111010"; -- Line 39   Column 14   Coefficient -0.02443695
         when "001001101110" => A <= "001001000110101001"; -- Line 39   Column 15   Coefficient 0.14224625
         when "001001101111" => A <= "001000110101000000"; -- Line 39   Column 16   Coefficient 0.13793945
         when "001001110000" => A <= "111111010000101110"; -- Line 40   Column 1   Coefficient -0.01154327
         when "001001110001" => A <= "000000001001011000"; -- Line 40   Column 2   Coefficient 0.00228882
         when "001001110010" => A <= "111111111111110100"; -- Line 40   Column 3   Coefficient -0.00004578
         when "001001110011" => A <= "000000000000000000"; -- Line 40   Column 4   Coefficient 0.00000000
         when "001001110100" => A <= "000000000000000000"; -- Line 40   Column 5   Coefficient 0.00000000
         when "001001110101" => A <= "000000000000000000"; -- Line 40   Column 6   Coefficient 0.00000000
         when "001001110110" => A <= "000000000000000000"; -- Line 40   Column 7   Coefficient 0.00000000
         when "001001110111" => A <= "000000000000000000"; -- Line 40   Column 8   Coefficient 0.00000000
         when "001001111000" => A <= "000000000000000000"; -- Line 40   Column 9   Coefficient 0.00000000
         when "001001111001" => A <= "000000000000000000"; -- Line 40   Column 10   Coefficient 0.00000000
         when "001001111010" => A <= "000000000000000000"; -- Line 40   Column 11   Coefficient 0.00000000
         when "001001111011" => A <= "000000000000000000"; -- Line 40   Column 12   Coefficient 0.00000000
         when "001001111100" => A <= "111111111111001011"; -- Line 40   Column 13   Coefficient -0.00020218
         when "001001111101" => A <= "111110100110010011"; -- Line 40   Column 14   Coefficient -0.02190018
         when "001001111110" => A <= "000111100110110001"; -- Line 40   Column 15   Coefficient 0.11883926
         when "001001111111" => A <= "001010011001111000"; -- Line 40   Column 16   Coefficient 0.16256714
         when "001010000000" => A <= "111110111010000001"; -- Line 41   Column 1   Coefficient -0.01708603
         when "001010000001" => A <= "000000010001001000"; -- Line 41   Column 2   Coefficient 0.00418091
         when "001010000010" => A <= "111111111111100110"; -- Line 41   Column 3   Coefficient -0.00009918
         when "001010000011" => A <= "000000000000000000"; -- Line 41   Column 4   Coefficient 0.00000000
         when "001010000100" => A <= "000000000000000000"; -- Line 41   Column 5   Coefficient 0.00000000
         when "001010000101" => A <= "000000000000000000"; -- Line 41   Column 6   Coefficient 0.00000000
         when "001010000110" => A <= "000000000000000000"; -- Line 41   Column 7   Coefficient 0.00000000
         when "001010000111" => A <= "000000000000000000"; -- Line 41   Column 8   Coefficient 0.00000000
         when "001010001000" => A <= "000000000000000000"; -- Line 41   Column 9   Coefficient 0.00000000
         when "001010001001" => A <= "000000000000000000"; -- Line 41   Column 10   Coefficient 0.00000000
         when "001010001010" => A <= "000000000000000000"; -- Line 41   Column 11   Coefficient 0.00000000
         when "001010001011" => A <= "000000000000000000"; -- Line 41   Column 12   Coefficient 0.00000000
         when "001010001100" => A <= "000000000000000011"; -- Line 41   Column 13   Coefficient 0.00001144
         when "001010001101" => A <= "111110110001100001"; -- Line 41   Column 14   Coefficient -0.01916122
         when "001010001110" => A <= "000110000101110011"; -- Line 41   Column 15   Coefficient 0.09516525
         when "001010001111" => A <= "001011111101111010"; -- Line 41   Column 16   Coefficient 0.18698883
         when "001010010000" => A <= "111110011010010101"; -- Line 42   Column 1   Coefficient -0.02482224
         when "001010010001" => A <= "000000011001110100"; -- Line 42   Column 2   Coefficient 0.00630188
         when "001010010010" => A <= "000000000000000111"; -- Line 42   Column 3   Coefficient 0.00002670
         when "001010010011" => A <= "000000000000000000"; -- Line 42   Column 4   Coefficient 0.00000000
         when "001010010100" => A <= "000000000000000000"; -- Line 42   Column 5   Coefficient 0.00000000
         when "001010010101" => A <= "000000000000000000"; -- Line 42   Column 6   Coefficient 0.00000000
         when "001010010110" => A <= "000000000000000000"; -- Line 42   Column 7   Coefficient 0.00000000
         when "001010010111" => A <= "000000000000000000"; -- Line 42   Column 8   Coefficient 0.00000000
         when "001010011000" => A <= "000000000000000000"; -- Line 42   Column 9   Coefficient 0.00000000
         when "001010011001" => A <= "000000000000000000"; -- Line 42   Column 10   Coefficient 0.00000000
         when "001010011010" => A <= "000000000000000000"; -- Line 42   Column 11   Coefficient 0.00000000
         when "001010011011" => A <= "000000000000000000"; -- Line 42   Column 12   Coefficient 0.00000000
         when "001010011100" => A <= "000000000000001001"; -- Line 42   Column 13   Coefficient 0.00003433
         when "001010011101" => A <= "111111000100111001"; -- Line 42   Column 14   Coefficient -0.01443100
         when "001010011110" => A <= "000100010010000101"; -- Line 42   Column 15   Coefficient 0.06691360
         when "001010011111" => A <= "001101110100101001"; -- Line 42   Column 16   Coefficient 0.21597672
         when "001010100000" => A <= "111101111110110001"; -- Line 43   Column 1   Coefficient -0.03155136
         when "001010100001" => A <= "000000100001110011"; -- Line 43   Column 2   Coefficient 0.00825119
         when "001010100010" => A <= "000000000000110011"; -- Line 43   Column 3   Coefficient 0.00019455
         when "001010100011" => A <= "000000000000000000"; -- Line 43   Column 4   Coefficient 0.00000000
         when "001010100100" => A <= "000000000000000000"; -- Line 43   Column 5   Coefficient 0.00000000
         when "001010100101" => A <= "000000000000000000"; -- Line 43   Column 6   Coefficient 0.00000000
         when "001010100110" => A <= "000000000000000000"; -- Line 43   Column 7   Coefficient 0.00000000
         when "001010100111" => A <= "000000000000000000"; -- Line 43   Column 8   Coefficient 0.00000000
         when "001010101000" => A <= "000000000000000000"; -- Line 43   Column 9   Coefficient 0.00000000
         when "001010101001" => A <= "000000000000000000"; -- Line 43   Column 10   Coefficient 0.00000000
         when "001010101010" => A <= "000000000000000000"; -- Line 43   Column 11   Coefficient 0.00000000
         when "001010101011" => A <= "000000000000000000"; -- Line 43   Column 12   Coefficient 0.00000000
         when "001010101100" => A <= "000000000000000000"; -- Line 43   Column 13   Coefficient 0.00000000
         when "001010101101" => A <= "111111011001111001"; -- Line 43   Column 14   Coefficient -0.00930405
         when "001010101110" => A <= "000010011110111100"; -- Line 43   Column 15   Coefficient 0.03880310
         when "001010101111" => A <= "001111100101110011"; -- Line 43   Column 16   Coefficient 0.24360275
         when "001010110000" => A <= "111101011101101101"; -- Line 44   Column 1   Coefficient -0.03962326
         when "001010110001" => A <= "000000101011110101"; -- Line 44   Column 2   Coefficient 0.01070023
         when "001010110010" => A <= "000000000001100101"; -- Line 44   Column 3   Coefficient 0.00038528
         when "001010110011" => A <= "000000000000000000"; -- Line 44   Column 4   Coefficient 0.00000000
         when "001010110100" => A <= "000000000000000000"; -- Line 44   Column 5   Coefficient 0.00000000
         when "001010110101" => A <= "000000000000000000"; -- Line 44   Column 6   Coefficient 0.00000000
         when "001010110110" => A <= "000000000000000000"; -- Line 44   Column 7   Coefficient 0.00000000
         when "001010110111" => A <= "000000000000000000"; -- Line 44   Column 8   Coefficient 0.00000000
         when "001010111000" => A <= "000000000000000000"; -- Line 44   Column 9   Coefficient 0.00000000
         when "001010111001" => A <= "000000000000000000"; -- Line 44   Column 10   Coefficient 0.00000000
         when "001010111010" => A <= "000000000000000000"; -- Line 44   Column 11   Coefficient 0.00000000
         when "001010111011" => A <= "000000000000000000"; -- Line 44   Column 12   Coefficient 0.00000000
         when "001010111100" => A <= "000000000000000000"; -- Line 44   Column 13   Coefficient 0.00000000
         when "001010111101" => A <= "111111110001010101"; -- Line 44   Column 14   Coefficient -0.00358200
         when "001010111110" => A <= "000000100101011001"; -- Line 44   Column 15   Coefficient 0.00912857
         when "001010111111" => A <= "010001011110001011"; -- Line 44   Column 16   Coefficient 0.27299118
         when "001011000000" => A <= "111101000110110001"; -- Line 45   Column 1   Coefficient -0.04522324
         when "001011000001" => A <= "000000110100010110"; -- Line 45   Column 2   Coefficient 0.01277924
         when "001011000010" => A <= "000000000010010101"; -- Line 45   Column 3   Coefficient 0.00056839
         when "001011000011" => A <= "000000000000000000"; -- Line 45   Column 4   Coefficient 0.00000000
         when "001011000100" => A <= "000000000000000000"; -- Line 45   Column 5   Coefficient 0.00000000
         when "001011000101" => A <= "000000000000000000"; -- Line 45   Column 6   Coefficient 0.00000000
         when "001011000110" => A <= "000000000000000000"; -- Line 45   Column 7   Coefficient 0.00000000
         when "001011000111" => A <= "000000000000000000"; -- Line 45   Column 8   Coefficient 0.00000000
         when "001011001000" => A <= "000000000000000000"; -- Line 45   Column 9   Coefficient 0.00000000
         when "001011001001" => A <= "000000000000000000"; -- Line 45   Column 10   Coefficient 0.00000000
         when "001011001010" => A <= "000000000000000000"; -- Line 45   Column 11   Coefficient 0.00000000
         when "001011001011" => A <= "000000000000000000"; -- Line 45   Column 12   Coefficient 0.00000000
         when "001011001100" => A <= "000000000000000000"; -- Line 45   Column 13   Coefficient 0.00000000
         when "001011001101" => A <= "000000000111011010"; -- Line 45   Column 14   Coefficient 0.00180817
         when "001011001110" => A <= "111110110101100100"; -- Line 45   Column 15   Coefficient -0.01817322
         when "001011001111" => A <= "010011000101100111"; -- Line 45   Column 16   Coefficient 0.29824448
         when "001011010000" => A <= "111101100111001110"; -- Line 46   Column 1   Coefficient -0.03730011
         when "001011010001" => A <= "000000110010101110"; -- Line 46   Column 2   Coefficient 0.01238251
         when "001011010010" => A <= "000000000001111110"; -- Line 46   Column 3   Coefficient 0.00048065
         when "001011010011" => A <= "000000000000000000"; -- Line 46   Column 4   Coefficient 0.00000000
         when "001011010100" => A <= "000000000000000000"; -- Line 46   Column 5   Coefficient 0.00000000
         when "001011010101" => A <= "000000000000000000"; -- Line 46   Column 6   Coefficient 0.00000000
         when "001011010110" => A <= "000000000000000000"; -- Line 46   Column 7   Coefficient 0.00000000
         when "001011010111" => A <= "000000000000000000"; -- Line 46   Column 8   Coefficient 0.00000000
         when "001011011000" => A <= "000000000000000000"; -- Line 46   Column 9   Coefficient 0.00000000
         when "001011011001" => A <= "000000000000000000"; -- Line 46   Column 10   Coefficient 0.00000000
         when "001011011010" => A <= "000000000000000000"; -- Line 46   Column 11   Coefficient 0.00000000
         when "001011011011" => A <= "000000000000000000"; -- Line 46   Column 12   Coefficient 0.00000000
         when "001011011100" => A <= "000000000000000000"; -- Line 46   Column 13   Coefficient 0.00000000
         when "001011011101" => A <= "000000001111000010"; -- Line 46   Column 14   Coefficient 0.00366974
         when "001011011110" => A <= "111110000010011110"; -- Line 46   Column 15   Coefficient -0.03064728
         when "001011011111" => A <= "010011010010100110"; -- Line 46   Column 16   Coefficient 0.30141449
         when "001011100000" => A <= "111110100000101100"; -- Line 47   Column 1   Coefficient -0.02326965
         when "001011100001" => A <= "000000101101010111"; -- Line 47   Column 2   Coefficient 0.01107407
         when "001011100010" => A <= "000000000001000010"; -- Line 47   Column 3   Coefficient 0.00025177
         when "001011100011" => A <= "000000000000000000"; -- Line 47   Column 4   Coefficient 0.00000000
         when "001011100100" => A <= "000000000000000000"; -- Line 47   Column 5   Coefficient 0.00000000
         when "001011100101" => A <= "000000000000000000"; -- Line 47   Column 6   Coefficient 0.00000000
         when "001011100110" => A <= "000000000000000000"; -- Line 47   Column 7   Coefficient 0.00000000
         when "001011100111" => A <= "000000000000000000"; -- Line 47   Column 8   Coefficient 0.00000000
         when "001011101000" => A <= "000000000000000000"; -- Line 47   Column 9   Coefficient 0.00000000
         when "001011101001" => A <= "000000000000000000"; -- Line 47   Column 10   Coefficient 0.00000000
         when "001011101010" => A <= "000000000000000000"; -- Line 47   Column 11   Coefficient 0.00000000
         when "001011101011" => A <= "000000000000000000"; -- Line 47   Column 12   Coefficient 0.00000000
         when "001011101100" => A <= "000000000000000000"; -- Line 47   Column 13   Coefficient 0.00000000
         when "001011101101" => A <= "000000010000011000"; -- Line 47   Column 14   Coefficient 0.00399780
         when "001011101110" => A <= "111101101011101110"; -- Line 47   Column 15   Coefficient -0.03620148
         when "001011101111" => A <= "010010110100110100"; -- Line 47   Column 16   Coefficient 0.29414368
         when "001011110000" => A <= "111111101010001000"; -- Line 48   Column 1   Coefficient -0.00534058
         when "001011110001" => A <= "000000100010100100"; -- Line 48   Column 2   Coefficient 0.00843811
         when "001011110010" => A <= "000000000001001000"; -- Line 48   Column 3   Coefficient 0.00027466
         when "001011110011" => A <= "000000000000000000"; -- Line 48   Column 4   Coefficient 0.00000000
         when "001011110100" => A <= "000000000000000000"; -- Line 48   Column 5   Coefficient 0.00000000
         when "001011110101" => A <= "000000000000000000"; -- Line 48   Column 6   Coefficient 0.00000000
         when "001011110110" => A <= "000000000000000000"; -- Line 48   Column 7   Coefficient 0.00000000
         when "001011110111" => A <= "000000000000000000"; -- Line 48   Column 8   Coefficient 0.00000000
         when "001011111000" => A <= "000000000000000000"; -- Line 48   Column 9   Coefficient 0.00000000
         when "001011111001" => A <= "000000000000000000"; -- Line 48   Column 10   Coefficient 0.00000000
         when "001011111010" => A <= "000000000000000000"; -- Line 48   Column 11   Coefficient 0.00000000
         when "001011111011" => A <= "000000000000000000"; -- Line 48   Column 12   Coefficient 0.00000000
         when "001011111100" => A <= "000000000000000000"; -- Line 48   Column 13   Coefficient 0.00000000
         when "001011111101" => A <= "000000001111111100"; -- Line 48   Column 14   Coefficient 0.00389099
         when "001011111110" => A <= "111101100000101101"; -- Line 48   Column 15   Coefficient -0.03889084
         when "001011111111" => A <= "010010000001100011"; -- Line 48   Column 16   Coefficient 0.28162766
         when "001100000000" => A <= "000000111110100110"; -- Line 49   Column 1   Coefficient 0.01528168
         when "001100000001" => A <= "000000010110010000"; -- Line 49   Column 2   Coefficient 0.00543213
         when "001100000010" => A <= "000000000001001011"; -- Line 49   Column 3   Coefficient 0.00028610
         when "001100000011" => A <= "000000000000000000"; -- Line 49   Column 4   Coefficient 0.00000000
         when "001100000100" => A <= "000000000000000000"; -- Line 49   Column 5   Coefficient 0.00000000
         when "001100000101" => A <= "000000000000000000"; -- Line 49   Column 6   Coefficient 0.00000000
         when "001100000110" => A <= "000000000000000000"; -- Line 49   Column 7   Coefficient 0.00000000
         when "001100000111" => A <= "000000000000000000"; -- Line 49   Column 8   Coefficient 0.00000000
         when "001100001000" => A <= "000000000000000000"; -- Line 49   Column 9   Coefficient 0.00000000
         when "001100001001" => A <= "000000000000000000"; -- Line 49   Column 10   Coefficient 0.00000000
         when "001100001010" => A <= "000000000000000000"; -- Line 49   Column 11   Coefficient 0.00000000
         when "001100001011" => A <= "000000000000000000"; -- Line 49   Column 12   Coefficient 0.00000000
         when "001100001100" => A <= "000000000000000000"; -- Line 49   Column 13   Coefficient 0.00000000
         when "001100001101" => A <= "000000001101001100"; -- Line 49   Column 14   Coefficient 0.00321960
         when "001100001110" => A <= "111101100010001110"; -- Line 49   Column 15   Coefficient -0.03852081
         when "001100001111" => A <= "010000111010100101"; -- Line 49   Column 16   Coefficient 0.26430130
         when "001100010000" => A <= "000010000100001011"; -- Line 50   Column 1   Coefficient 0.03226852
         when "001100010001" => A <= "000000010100110111"; -- Line 50   Column 2   Coefficient 0.00509262
         when "001100010010" => A <= "111111111110110111"; -- Line 50   Column 3   Coefficient -0.00027847
         when "001100010011" => A <= "000000000000000000"; -- Line 50   Column 4   Coefficient 0.00000000
         when "001100010100" => A <= "000000000000000000"; -- Line 50   Column 5   Coefficient 0.00000000
         when "001100010101" => A <= "000000000000000000"; -- Line 50   Column 6   Coefficient 0.00000000
         when "001100010110" => A <= "000000000000000000"; -- Line 50   Column 7   Coefficient 0.00000000
         when "001100010111" => A <= "000000000000000000"; -- Line 50   Column 8   Coefficient 0.00000000
         when "001100011000" => A <= "000000000000000000"; -- Line 50   Column 9   Coefficient 0.00000000
         when "001100011001" => A <= "000000000000000000"; -- Line 50   Column 10   Coefficient 0.00000000
         when "001100011010" => A <= "000000000000000000"; -- Line 50   Column 11   Coefficient 0.00000000
         when "001100011011" => A <= "000000000000000000"; -- Line 50   Column 12   Coefficient 0.00000000
         when "001100011100" => A <= "000000000000000000"; -- Line 50   Column 13   Coefficient 0.00000000
         when "001100011101" => A <= "000000001010110110"; -- Line 50   Column 14   Coefficient 0.00264740
         when "001100011110" => A <= "111101100010101111"; -- Line 50   Column 15   Coefficient -0.03839493
         when "001100011111" => A <= "001111111010100001"; -- Line 50   Column 16   Coefficient 0.24866104
         when "001100100000" => A <= "000011001010010011"; -- Line 51   Column 1   Coefficient 0.04938889
         when "001100100001" => A <= "000000010100111001"; -- Line 51   Column 2   Coefficient 0.00510025
         when "001100100010" => A <= "111111111100011110"; -- Line 51   Column 3   Coefficient -0.00086212
         when "001100100011" => A <= "111111111111111111"; -- Line 51   Column 4   Coefficient -0.00000381
         when "001100100100" => A <= "000000000000000000"; -- Line 51   Column 5   Coefficient 0.00000000
         when "001100100101" => A <= "000000000000000000"; -- Line 51   Column 6   Coefficient 0.00000000
         when "001100100110" => A <= "000000000000000000"; -- Line 51   Column 7   Coefficient 0.00000000
         when "001100100111" => A <= "000000000000000000"; -- Line 51   Column 8   Coefficient 0.00000000
         when "001100101000" => A <= "000000000000000000"; -- Line 51   Column 9   Coefficient 0.00000000
         when "001100101001" => A <= "000000000000000000"; -- Line 51   Column 10   Coefficient 0.00000000
         when "001100101010" => A <= "000000000000000000"; -- Line 51   Column 11   Coefficient 0.00000000
         when "001100101011" => A <= "000000000000000000"; -- Line 51   Column 12   Coefficient 0.00000000
         when "001100101100" => A <= "000000000000000000"; -- Line 51   Column 13   Coefficient 0.00000000
         when "001100101101" => A <= "000000001000010011"; -- Line 51   Column 14   Coefficient 0.00202560
         when "001100101110" => A <= "111101100110110000"; -- Line 51   Column 15   Coefficient -0.03741455
         when "001100101111" => A <= "001110110101010100"; -- Line 51   Column 16   Coefficient 0.23176575
         when "001100110000" => A <= "000100010011001101"; -- Line 52   Column 1   Coefficient 0.06718826
         when "001100110001" => A <= "000000010111101010"; -- Line 52   Column 2   Coefficient 0.00577545
         when "001100110010" => A <= "111111111001000110"; -- Line 52   Column 3   Coefficient -0.00168610
         when "001100110011" => A <= "000000000000000011"; -- Line 52   Column 4   Coefficient 0.00001144
         when "001100110100" => A <= "000000000000000000"; -- Line 52   Column 5   Coefficient 0.00000000
         when "001100110101" => A <= "000000000000000000"; -- Line 52   Column 6   Coefficient 0.00000000
         when "001100110110" => A <= "000000000000000000"; -- Line 52   Column 7   Coefficient 0.00000000
         when "001100110111" => A <= "000000000000000000"; -- Line 52   Column 8   Coefficient 0.00000000
         when "001100111000" => A <= "000000000000000000"; -- Line 52   Column 9   Coefficient 0.00000000
         when "001100111001" => A <= "000000000000000000"; -- Line 52   Column 10   Coefficient 0.00000000
         when "001100111010" => A <= "000000000000000000"; -- Line 52   Column 11   Coefficient 0.00000000
         when "001100111011" => A <= "000000000000000000"; -- Line 52   Column 12   Coefficient 0.00000000
         when "001100111100" => A <= "000000000000000000"; -- Line 52   Column 13   Coefficient 0.00000000
         when "001100111101" => A <= "000000000011111000"; -- Line 52   Column 14   Coefficient 0.00094604
         when "001100111110" => A <= "111101110100001010"; -- Line 52   Column 15   Coefficient -0.03414154
         when "001100111111" => A <= "001101100011111111"; -- Line 52   Column 16   Coefficient 0.21191025
         when "001101000000" => A <= "000101100000010101"; -- Line 53   Column 1   Coefficient 0.08601761
         when "001101000001" => A <= "000000011000110111"; -- Line 53   Column 2   Coefficient 0.00606918
         when "001101000010" => A <= "111111110110011111"; -- Line 53   Column 3   Coefficient -0.00232315
         when "001101000011" => A <= "000000000000000110"; -- Line 53   Column 4   Coefficient 0.00002289
         when "001101000100" => A <= "000000000000000000"; -- Line 53   Column 5   Coefficient 0.00000000
         when "001101000101" => A <= "000000000000000000"; -- Line 53   Column 6   Coefficient 0.00000000
         when "001101000110" => A <= "000000000000000000"; -- Line 53   Column 7   Coefficient 0.00000000
         when "001101000111" => A <= "000000000000000000"; -- Line 53   Column 8   Coefficient 0.00000000
         when "001101001000" => A <= "000000000000000000"; -- Line 53   Column 9   Coefficient 0.00000000
         when "001101001001" => A <= "000000000000000000"; -- Line 53   Column 10   Coefficient 0.00000000
         when "001101001010" => A <= "000000000000000000"; -- Line 53   Column 11   Coefficient 0.00000000
         when "001101001011" => A <= "000000000000000000"; -- Line 53   Column 12   Coefficient 0.00000000
         when "001101001100" => A <= "000000000000000000"; -- Line 53   Column 13   Coefficient 0.00000000
         when "001101001101" => A <= "111111111111010011"; -- Line 53   Column 14   Coefficient -0.00017166
         when "001101001110" => A <= "111110000101010011"; -- Line 53   Column 15   Coefficient -0.02995682
         when "001101001111" => A <= "001100001011101000"; -- Line 53   Column 16   Coefficient 0.19033813
         when "001101010000" => A <= "000111000101010101"; -- Line 54   Column 1   Coefficient 0.11067581
         when "001101010001" => A <= "000000000100100100"; -- Line 54   Column 2   Coefficient 0.00111389
         when "001101010010" => A <= "111111111010111001"; -- Line 54   Column 3   Coefficient -0.00124741
         when "001101010011" => A <= "000000000000000100"; -- Line 54   Column 4   Coefficient 0.00001526
         when "001101010100" => A <= "000000000000000000"; -- Line 54   Column 5   Coefficient 0.00000000
         when "001101010101" => A <= "000000000000000000"; -- Line 54   Column 6   Coefficient 0.00000000
         when "001101010110" => A <= "000000000000000000"; -- Line 54   Column 7   Coefficient 0.00000000
         when "001101010111" => A <= "000000000000000000"; -- Line 54   Column 8   Coefficient 0.00000000
         when "001101011000" => A <= "000000000000000000"; -- Line 54   Column 9   Coefficient 0.00000000
         when "001101011001" => A <= "000000000000000000"; -- Line 54   Column 10   Coefficient 0.00000000
         when "001101011010" => A <= "000000000000000000"; -- Line 54   Column 11   Coefficient 0.00000000
         when "001101011011" => A <= "000000000000000000"; -- Line 54   Column 12   Coefficient 0.00000000
         when "001101011100" => A <= "000000000000000000"; -- Line 54   Column 13   Coefficient 0.00000000
         when "001101011101" => A <= "111111111110010010"; -- Line 54   Column 14   Coefficient -0.00041962
         when "001101011110" => A <= "111110010000110000"; -- Line 54   Column 15   Coefficient -0.02716064
         when "001101011111" => A <= "001010101100000111"; -- Line 54   Column 16   Coefficient 0.16701889
         when "001101100000" => A <= "001000110101000000"; -- Line 55   Column 1   Coefficient 0.13793945
         when "001101100001" => A <= "111111100111100010"; -- Line 55   Column 2   Coefficient -0.00597382
         when "001101100010" => A <= "000000000010010011"; -- Line 55   Column 3   Coefficient 0.00056076
         when "001101100011" => A <= "000000000000000011"; -- Line 55   Column 4   Coefficient 0.00001144
         when "001101100100" => A <= "000000000000000000"; -- Line 55   Column 5   Coefficient 0.00000000
         when "001101100101" => A <= "000000000000000000"; -- Line 55   Column 6   Coefficient 0.00000000
         when "001101100110" => A <= "000000000000000000"; -- Line 55   Column 7   Coefficient 0.00000000
         when "001101100111" => A <= "000000000000000000"; -- Line 55   Column 8   Coefficient 0.00000000
         when "001101101000" => A <= "000000000000000000"; -- Line 55   Column 9   Coefficient 0.00000000
         when "001101101001" => A <= "000000000000000000"; -- Line 55   Column 10   Coefficient 0.00000000
         when "001101101010" => A <= "000000000000000000"; -- Line 55   Column 11   Coefficient 0.00000000
         when "001101101011" => A <= "000000000000000000"; -- Line 55   Column 12   Coefficient 0.00000000
         when "001101101100" => A <= "000000000000000000"; -- Line 55   Column 13   Coefficient 0.00000000
         when "001101101101" => A <= "111111111110100110"; -- Line 55   Column 14   Coefficient -0.00034332
         when "001101101110" => A <= "111110011011111010"; -- Line 55   Column 15   Coefficient -0.02443695
         when "001101101111" => A <= "001001000110101001"; -- Line 55   Column 16   Coefficient 0.14224625
         when "001101110000" => A <= "001010011001111000"; -- Line 56   Column 1   Coefficient 0.16256714
         when "001101110001" => A <= "111111010000101110"; -- Line 56   Column 2   Coefficient -0.01154327
         when "001101110010" => A <= "000000001001011000"; -- Line 56   Column 3   Coefficient 0.00228882
         when "001101110011" => A <= "111111111111110100"; -- Line 56   Column 4   Coefficient -0.00004578
         when "001101110100" => A <= "000000000000000000"; -- Line 56   Column 5   Coefficient 0.00000000
         when "001101110101" => A <= "000000000000000000"; -- Line 56   Column 6   Coefficient 0.00000000
         when "001101110110" => A <= "000000000000000000"; -- Line 56   Column 7   Coefficient 0.00000000
         when "001101110111" => A <= "000000000000000000"; -- Line 56   Column 8   Coefficient 0.00000000
         when "001101111000" => A <= "000000000000000000"; -- Line 56   Column 9   Coefficient 0.00000000
         when "001101111001" => A <= "000000000000000000"; -- Line 56   Column 10   Coefficient 0.00000000
         when "001101111010" => A <= "000000000000000000"; -- Line 56   Column 11   Coefficient 0.00000000
         when "001101111011" => A <= "000000000000000000"; -- Line 56   Column 12   Coefficient 0.00000000
         when "001101111100" => A <= "000000000000000000"; -- Line 56   Column 13   Coefficient 0.00000000
         when "001101111101" => A <= "111111111111001011"; -- Line 56   Column 14   Coefficient -0.00020218
         when "001101111110" => A <= "111110100110010011"; -- Line 56   Column 15   Coefficient -0.02190018
         when "001101111111" => A <= "000111100110110001"; -- Line 56   Column 16   Coefficient 0.11883926
         when "001110000000" => A <= "001011111101111010"; -- Line 57   Column 1   Coefficient 0.18698883
         when "001110000001" => A <= "111110111010000001"; -- Line 57   Column 2   Coefficient -0.01708603
         when "001110000010" => A <= "000000010001001000"; -- Line 57   Column 3   Coefficient 0.00418091
         when "001110000011" => A <= "111111111111100110"; -- Line 57   Column 4   Coefficient -0.00009918
         when "001110000100" => A <= "000000000000000000"; -- Line 57   Column 5   Coefficient 0.00000000
         when "001110000101" => A <= "000000000000000000"; -- Line 57   Column 6   Coefficient 0.00000000
         when "001110000110" => A <= "000000000000000000"; -- Line 57   Column 7   Coefficient 0.00000000
         when "001110000111" => A <= "000000000000000000"; -- Line 57   Column 8   Coefficient 0.00000000
         when "001110001000" => A <= "000000000000000000"; -- Line 57   Column 9   Coefficient 0.00000000
         when "001110001001" => A <= "000000000000000000"; -- Line 57   Column 10   Coefficient 0.00000000
         when "001110001010" => A <= "000000000000000000"; -- Line 57   Column 11   Coefficient 0.00000000
         when "001110001011" => A <= "000000000000000000"; -- Line 57   Column 12   Coefficient 0.00000000
         when "001110001100" => A <= "000000000000000000"; -- Line 57   Column 13   Coefficient 0.00000000
         when "001110001101" => A <= "000000000000000011"; -- Line 57   Column 14   Coefficient 0.00001144
         when "001110001110" => A <= "111110110001100001"; -- Line 57   Column 15   Coefficient -0.01916122
         when "001110001111" => A <= "000110000101110011"; -- Line 57   Column 16   Coefficient 0.09516525
         when "001110010000" => A <= "001101110100101001"; -- Line 58   Column 1   Coefficient 0.21597672
         when "001110010001" => A <= "111110011010010101"; -- Line 58   Column 2   Coefficient -0.02482224
         when "001110010010" => A <= "000000011001110100"; -- Line 58   Column 3   Coefficient 0.00630188
         when "001110010011" => A <= "000000000000000111"; -- Line 58   Column 4   Coefficient 0.00002670
         when "001110010100" => A <= "000000000000000000"; -- Line 58   Column 5   Coefficient 0.00000000
         when "001110010101" => A <= "000000000000000000"; -- Line 58   Column 6   Coefficient 0.00000000
         when "001110010110" => A <= "000000000000000000"; -- Line 58   Column 7   Coefficient 0.00000000
         when "001110010111" => A <= "000000000000000000"; -- Line 58   Column 8   Coefficient 0.00000000
         when "001110011000" => A <= "000000000000000000"; -- Line 58   Column 9   Coefficient 0.00000000
         when "001110011001" => A <= "000000000000000000"; -- Line 58   Column 10   Coefficient 0.00000000
         when "001110011010" => A <= "000000000000000000"; -- Line 58   Column 11   Coefficient 0.00000000
         when "001110011011" => A <= "000000000000000000"; -- Line 58   Column 12   Coefficient 0.00000000
         when "001110011100" => A <= "000000000000000000"; -- Line 58   Column 13   Coefficient 0.00000000
         when "001110011101" => A <= "000000000000001001"; -- Line 58   Column 14   Coefficient 0.00003433
         when "001110011110" => A <= "111111000100111001"; -- Line 58   Column 15   Coefficient -0.01443100
         when "001110011111" => A <= "000100010010000101"; -- Line 58   Column 16   Coefficient 0.06691360
         when "001110100000" => A <= "001111100101110011"; -- Line 59   Column 1   Coefficient 0.24360275
         when "001110100001" => A <= "111101111110110001"; -- Line 59   Column 2   Coefficient -0.03155136
         when "001110100010" => A <= "000000100001110011"; -- Line 59   Column 3   Coefficient 0.00825119
         when "001110100011" => A <= "000000000000110011"; -- Line 59   Column 4   Coefficient 0.00019455
         when "001110100100" => A <= "000000000000000000"; -- Line 59   Column 5   Coefficient 0.00000000
         when "001110100101" => A <= "000000000000000000"; -- Line 59   Column 6   Coefficient 0.00000000
         when "001110100110" => A <= "000000000000000000"; -- Line 59   Column 7   Coefficient 0.00000000
         when "001110100111" => A <= "000000000000000000"; -- Line 59   Column 8   Coefficient 0.00000000
         when "001110101000" => A <= "000000000000000000"; -- Line 59   Column 9   Coefficient 0.00000000
         when "001110101001" => A <= "000000000000000000"; -- Line 59   Column 10   Coefficient 0.00000000
         when "001110101010" => A <= "000000000000000000"; -- Line 59   Column 11   Coefficient 0.00000000
         when "001110101011" => A <= "000000000000000000"; -- Line 59   Column 12   Coefficient 0.00000000
         when "001110101100" => A <= "000000000000000000"; -- Line 59   Column 13   Coefficient 0.00000000
         when "001110101101" => A <= "000000000000000000"; -- Line 59   Column 14   Coefficient 0.00000000
         when "001110101110" => A <= "111111011001111001"; -- Line 59   Column 15   Coefficient -0.00930405
         when "001110101111" => A <= "000010011110111100"; -- Line 59   Column 16   Coefficient 0.03880310
         when "001110110000" => A <= "010001011110001011"; -- Line 60   Column 1   Coefficient 0.27299118
         when "001110110001" => A <= "111101011101101101"; -- Line 60   Column 2   Coefficient -0.03962326
         when "001110110010" => A <= "000000101011110101"; -- Line 60   Column 3   Coefficient 0.01070023
         when "001110110011" => A <= "000000000001100101"; -- Line 60   Column 4   Coefficient 0.00038528
         when "001110110100" => A <= "000000000000000000"; -- Line 60   Column 5   Coefficient 0.00000000
         when "001110110101" => A <= "000000000000000000"; -- Line 60   Column 6   Coefficient 0.00000000
         when "001110110110" => A <= "000000000000000000"; -- Line 60   Column 7   Coefficient 0.00000000
         when "001110110111" => A <= "000000000000000000"; -- Line 60   Column 8   Coefficient 0.00000000
         when "001110111000" => A <= "000000000000000000"; -- Line 60   Column 9   Coefficient 0.00000000
         when "001110111001" => A <= "000000000000000000"; -- Line 60   Column 10   Coefficient 0.00000000
         when "001110111010" => A <= "000000000000000000"; -- Line 60   Column 11   Coefficient 0.00000000
         when "001110111011" => A <= "000000000000000000"; -- Line 60   Column 12   Coefficient 0.00000000
         when "001110111100" => A <= "000000000000000000"; -- Line 60   Column 13   Coefficient 0.00000000
         when "001110111101" => A <= "000000000000000000"; -- Line 60   Column 14   Coefficient 0.00000000
         when "001110111110" => A <= "111111110001010101"; -- Line 60   Column 15   Coefficient -0.00358200
         when "001110111111" => A <= "000000100101011001"; -- Line 60   Column 16   Coefficient 0.00912857
         when "001111000000" => A <= "010011000101100111"; -- Line 61   Column 1   Coefficient 0.29824448
         when "001111000001" => A <= "111101000110110001"; -- Line 61   Column 2   Coefficient -0.04522324
         when "001111000010" => A <= "000000110100010110"; -- Line 61   Column 3   Coefficient 0.01277924
         when "001111000011" => A <= "000000000010010101"; -- Line 61   Column 4   Coefficient 0.00056839
         when "001111000100" => A <= "000000000000000000"; -- Line 61   Column 5   Coefficient 0.00000000
         when "001111000101" => A <= "000000000000000000"; -- Line 61   Column 6   Coefficient 0.00000000
         when "001111000110" => A <= "000000000000000000"; -- Line 61   Column 7   Coefficient 0.00000000
         when "001111000111" => A <= "000000000000000000"; -- Line 61   Column 8   Coefficient 0.00000000
         when "001111001000" => A <= "000000000000000000"; -- Line 61   Column 9   Coefficient 0.00000000
         when "001111001001" => A <= "000000000000000000"; -- Line 61   Column 10   Coefficient 0.00000000
         when "001111001010" => A <= "000000000000000000"; -- Line 61   Column 11   Coefficient 0.00000000
         when "001111001011" => A <= "000000000000000000"; -- Line 61   Column 12   Coefficient 0.00000000
         when "001111001100" => A <= "000000000000000000"; -- Line 61   Column 13   Coefficient 0.00000000
         when "001111001101" => A <= "000000000000000000"; -- Line 61   Column 14   Coefficient 0.00000000
         when "001111001110" => A <= "000000000111011010"; -- Line 61   Column 15   Coefficient 0.00180817
         when "001111001111" => A <= "111110110101100100"; -- Line 61   Column 16   Coefficient -0.01817322
         when "001111010000" => A <= "010011010010100110"; -- Line 62   Column 1   Coefficient 0.30141449
         when "001111010001" => A <= "111101100111001110"; -- Line 62   Column 2   Coefficient -0.03730011
         when "001111010010" => A <= "000000110010101110"; -- Line 62   Column 3   Coefficient 0.01238251
         when "001111010011" => A <= "000000000001111110"; -- Line 62   Column 4   Coefficient 0.00048065
         when "001111010100" => A <= "000000000000000000"; -- Line 62   Column 5   Coefficient 0.00000000
         when "001111010101" => A <= "000000000000000000"; -- Line 62   Column 6   Coefficient 0.00000000
         when "001111010110" => A <= "000000000000000000"; -- Line 62   Column 7   Coefficient 0.00000000
         when "001111010111" => A <= "000000000000000000"; -- Line 62   Column 8   Coefficient 0.00000000
         when "001111011000" => A <= "000000000000000000"; -- Line 62   Column 9   Coefficient 0.00000000
         when "001111011001" => A <= "000000000000000000"; -- Line 62   Column 10   Coefficient 0.00000000
         when "001111011010" => A <= "000000000000000000"; -- Line 62   Column 11   Coefficient 0.00000000
         when "001111011011" => A <= "000000000000000000"; -- Line 62   Column 12   Coefficient 0.00000000
         when "001111011100" => A <= "000000000000000000"; -- Line 62   Column 13   Coefficient 0.00000000
         when "001111011101" => A <= "000000000000000000"; -- Line 62   Column 14   Coefficient 0.00000000
         when "001111011110" => A <= "000000001111000010"; -- Line 62   Column 15   Coefficient 0.00366974
         when "001111011111" => A <= "111110000010011110"; -- Line 62   Column 16   Coefficient -0.03064728
         when "001111100000" => A <= "010010110100110100"; -- Line 63   Column 1   Coefficient 0.29414368
         when "001111100001" => A <= "111110100000101100"; -- Line 63   Column 2   Coefficient -0.02326965
         when "001111100010" => A <= "000000101101010111"; -- Line 63   Column 3   Coefficient 0.01107407
         when "001111100011" => A <= "000000000001000010"; -- Line 63   Column 4   Coefficient 0.00025177
         when "001111100100" => A <= "000000000000000000"; -- Line 63   Column 5   Coefficient 0.00000000
         when "001111100101" => A <= "000000000000000000"; -- Line 63   Column 6   Coefficient 0.00000000
         when "001111100110" => A <= "000000000000000000"; -- Line 63   Column 7   Coefficient 0.00000000
         when "001111100111" => A <= "000000000000000000"; -- Line 63   Column 8   Coefficient 0.00000000
         when "001111101000" => A <= "000000000000000000"; -- Line 63   Column 9   Coefficient 0.00000000
         when "001111101001" => A <= "000000000000000000"; -- Line 63   Column 10   Coefficient 0.00000000
         when "001111101010" => A <= "000000000000000000"; -- Line 63   Column 11   Coefficient 0.00000000
         when "001111101011" => A <= "000000000000000000"; -- Line 63   Column 12   Coefficient 0.00000000
         when "001111101100" => A <= "000000000000000000"; -- Line 63   Column 13   Coefficient 0.00000000
         when "001111101101" => A <= "000000000000000000"; -- Line 63   Column 14   Coefficient 0.00000000
         when "001111101110" => A <= "000000010000011000"; -- Line 63   Column 15   Coefficient 0.00399780
         when "001111101111" => A <= "111101101011101110"; -- Line 63   Column 16   Coefficient -0.03620148
         when "001111110000" => A <= "010010000001100011"; -- Line 64   Column 1   Coefficient 0.28162766
         when "001111110001" => A <= "111111101010001000"; -- Line 64   Column 2   Coefficient -0.00534058
         when "001111110010" => A <= "000000100010100100"; -- Line 64   Column 3   Coefficient 0.00843811
         when "001111110011" => A <= "000000000001001000"; -- Line 64   Column 4   Coefficient 0.00027466
         when "001111110100" => A <= "000000000000000000"; -- Line 64   Column 5   Coefficient 0.00000000
         when "001111110101" => A <= "000000000000000000"; -- Line 64   Column 6   Coefficient 0.00000000
         when "001111110110" => A <= "000000000000000000"; -- Line 64   Column 7   Coefficient 0.00000000
         when "001111110111" => A <= "000000000000000000"; -- Line 64   Column 8   Coefficient 0.00000000
         when "001111111000" => A <= "000000000000000000"; -- Line 64   Column 9   Coefficient 0.00000000
         when "001111111001" => A <= "000000000000000000"; -- Line 64   Column 10   Coefficient 0.00000000
         when "001111111010" => A <= "000000000000000000"; -- Line 64   Column 11   Coefficient 0.00000000
         when "001111111011" => A <= "000000000000000000"; -- Line 64   Column 12   Coefficient 0.00000000
         when "001111111100" => A <= "000000000000000000"; -- Line 64   Column 13   Coefficient 0.00000000
         when "001111111101" => A <= "000000000000000000"; -- Line 64   Column 14   Coefficient 0.00000000
         when "001111111110" => A <= "000000001111111100"; -- Line 64   Column 15   Coefficient 0.00389099
         when "001111111111" => A <= "111101100000101101"; -- Line 64   Column 16   Coefficient -0.03889084
         when "010000000000" => A <= "010000111010100101"; -- Line 65   Column 1   Coefficient 0.26430130
         when "010000000001" => A <= "000000111110100110"; -- Line 65   Column 2   Coefficient 0.01528168
         when "010000000010" => A <= "000000010110010000"; -- Line 65   Column 3   Coefficient 0.00543213
         when "010000000011" => A <= "000000000001001011"; -- Line 65   Column 4   Coefficient 0.00028610
         when "010000000100" => A <= "000000000000000000"; -- Line 65   Column 5   Coefficient 0.00000000
         when "010000000101" => A <= "000000000000000000"; -- Line 65   Column 6   Coefficient 0.00000000
         when "010000000110" => A <= "000000000000000000"; -- Line 65   Column 7   Coefficient 0.00000000
         when "010000000111" => A <= "000000000000000000"; -- Line 65   Column 8   Coefficient 0.00000000
         when "010000001000" => A <= "000000000000000000"; -- Line 65   Column 9   Coefficient 0.00000000
         when "010000001001" => A <= "000000000000000000"; -- Line 65   Column 10   Coefficient 0.00000000
         when "010000001010" => A <= "000000000000000000"; -- Line 65   Column 11   Coefficient 0.00000000
         when "010000001011" => A <= "000000000000000000"; -- Line 65   Column 12   Coefficient 0.00000000
         when "010000001100" => A <= "000000000000000000"; -- Line 65   Column 13   Coefficient 0.00000000
         when "010000001101" => A <= "000000000000000000"; -- Line 65   Column 14   Coefficient 0.00000000
         when "010000001110" => A <= "000000001101001100"; -- Line 65   Column 15   Coefficient 0.00321960
         when "010000001111" => A <= "111101100010001110"; -- Line 65   Column 16   Coefficient -0.03852081
         when "010000010000" => A <= "001111111010100001"; -- Line 66   Column 1   Coefficient 0.24866104
         when "010000010001" => A <= "000010000100001011"; -- Line 66   Column 2   Coefficient 0.03226852
         when "010000010010" => A <= "000000010100110111"; -- Line 66   Column 3   Coefficient 0.00509262
         when "010000010011" => A <= "111111111110110111"; -- Line 66   Column 4   Coefficient -0.00027847
         when "010000010100" => A <= "000000000000000000"; -- Line 66   Column 5   Coefficient 0.00000000
         when "010000010101" => A <= "000000000000000000"; -- Line 66   Column 6   Coefficient 0.00000000
         when "010000010110" => A <= "000000000000000000"; -- Line 66   Column 7   Coefficient 0.00000000
         when "010000010111" => A <= "000000000000000000"; -- Line 66   Column 8   Coefficient 0.00000000
         when "010000011000" => A <= "000000000000000000"; -- Line 66   Column 9   Coefficient 0.00000000
         when "010000011001" => A <= "000000000000000000"; -- Line 66   Column 10   Coefficient 0.00000000
         when "010000011010" => A <= "000000000000000000"; -- Line 66   Column 11   Coefficient 0.00000000
         when "010000011011" => A <= "000000000000000000"; -- Line 66   Column 12   Coefficient 0.00000000
         when "010000011100" => A <= "000000000000000000"; -- Line 66   Column 13   Coefficient 0.00000000
         when "010000011101" => A <= "000000000000000000"; -- Line 66   Column 14   Coefficient 0.00000000
         when "010000011110" => A <= "000000001010110110"; -- Line 66   Column 15   Coefficient 0.00264740
         when "010000011111" => A <= "111101100010101111"; -- Line 66   Column 16   Coefficient -0.03839493
         when "010000100000" => A <= "001110110101010100"; -- Line 67   Column 1   Coefficient 0.23176575
         when "010000100001" => A <= "000011001010010011"; -- Line 67   Column 2   Coefficient 0.04938889
         when "010000100010" => A <= "000000010100111001"; -- Line 67   Column 3   Coefficient 0.00510025
         when "010000100011" => A <= "111111111100011110"; -- Line 67   Column 4   Coefficient -0.00086212
         when "010000100100" => A <= "111111111111111111"; -- Line 67   Column 5   Coefficient -0.00000381
         when "010000100101" => A <= "000000000000000000"; -- Line 67   Column 6   Coefficient 0.00000000
         when "010000100110" => A <= "000000000000000000"; -- Line 67   Column 7   Coefficient 0.00000000
         when "010000100111" => A <= "000000000000000000"; -- Line 67   Column 8   Coefficient 0.00000000
         when "010000101000" => A <= "000000000000000000"; -- Line 67   Column 9   Coefficient 0.00000000
         when "010000101001" => A <= "000000000000000000"; -- Line 67   Column 10   Coefficient 0.00000000
         when "010000101010" => A <= "000000000000000000"; -- Line 67   Column 11   Coefficient 0.00000000
         when "010000101011" => A <= "000000000000000000"; -- Line 67   Column 12   Coefficient 0.00000000
         when "010000101100" => A <= "000000000000000000"; -- Line 67   Column 13   Coefficient 0.00000000
         when "010000101101" => A <= "000000000000000000"; -- Line 67   Column 14   Coefficient 0.00000000
         when "010000101110" => A <= "000000001000010011"; -- Line 67   Column 15   Coefficient 0.00202560
         when "010000101111" => A <= "111101100110110000"; -- Line 67   Column 16   Coefficient -0.03741455
         when "010000110000" => A <= "001101100011111111"; -- Line 68   Column 1   Coefficient 0.21191025
         when "010000110001" => A <= "000100010011001101"; -- Line 68   Column 2   Coefficient 0.06718826
         when "010000110010" => A <= "000000010111101010"; -- Line 68   Column 3   Coefficient 0.00577545
         when "010000110011" => A <= "111111111001000110"; -- Line 68   Column 4   Coefficient -0.00168610
         when "010000110100" => A <= "000000000000000011"; -- Line 68   Column 5   Coefficient 0.00001144
         when "010000110101" => A <= "000000000000000000"; -- Line 68   Column 6   Coefficient 0.00000000
         when "010000110110" => A <= "000000000000000000"; -- Line 68   Column 7   Coefficient 0.00000000
         when "010000110111" => A <= "000000000000000000"; -- Line 68   Column 8   Coefficient 0.00000000
         when "010000111000" => A <= "000000000000000000"; -- Line 68   Column 9   Coefficient 0.00000000
         when "010000111001" => A <= "000000000000000000"; -- Line 68   Column 10   Coefficient 0.00000000
         when "010000111010" => A <= "000000000000000000"; -- Line 68   Column 11   Coefficient 0.00000000
         when "010000111011" => A <= "000000000000000000"; -- Line 68   Column 12   Coefficient 0.00000000
         when "010000111100" => A <= "000000000000000000"; -- Line 68   Column 13   Coefficient 0.00000000
         when "010000111101" => A <= "000000000000000000"; -- Line 68   Column 14   Coefficient 0.00000000
         when "010000111110" => A <= "000000000011111000"; -- Line 68   Column 15   Coefficient 0.00094604
         when "010000111111" => A <= "111101110100001010"; -- Line 68   Column 16   Coefficient -0.03414154
         when "010001000000" => A <= "001100001011101000"; -- Line 69   Column 1   Coefficient 0.19033813
         when "010001000001" => A <= "000101100000010101"; -- Line 69   Column 2   Coefficient 0.08601761
         when "010001000010" => A <= "000000011000110111"; -- Line 69   Column 3   Coefficient 0.00606918
         when "010001000011" => A <= "111111110110011111"; -- Line 69   Column 4   Coefficient -0.00232315
         when "010001000100" => A <= "000000000000000110"; -- Line 69   Column 5   Coefficient 0.00002289
         when "010001000101" => A <= "000000000000000000"; -- Line 69   Column 6   Coefficient 0.00000000
         when "010001000110" => A <= "000000000000000000"; -- Line 69   Column 7   Coefficient 0.00000000
         when "010001000111" => A <= "000000000000000000"; -- Line 69   Column 8   Coefficient 0.00000000
         when "010001001000" => A <= "000000000000000000"; -- Line 69   Column 9   Coefficient 0.00000000
         when "010001001001" => A <= "000000000000000000"; -- Line 69   Column 10   Coefficient 0.00000000
         when "010001001010" => A <= "000000000000000000"; -- Line 69   Column 11   Coefficient 0.00000000
         when "010001001011" => A <= "000000000000000000"; -- Line 69   Column 12   Coefficient 0.00000000
         when "010001001100" => A <= "000000000000000000"; -- Line 69   Column 13   Coefficient 0.00000000
         when "010001001101" => A <= "000000000000000000"; -- Line 69   Column 14   Coefficient 0.00000000
         when "010001001110" => A <= "111111111111010011"; -- Line 69   Column 15   Coefficient -0.00017166
         when "010001001111" => A <= "111110000101010011"; -- Line 69   Column 16   Coefficient -0.02995682
         when "010001010000" => A <= "001010101100000111"; -- Line 70   Column 1   Coefficient 0.16701889
         when "010001010001" => A <= "000111000101010101"; -- Line 70   Column 2   Coefficient 0.11067581
         when "010001010010" => A <= "000000000100100100"; -- Line 70   Column 3   Coefficient 0.00111389
         when "010001010011" => A <= "111111111010111001"; -- Line 70   Column 4   Coefficient -0.00124741
         when "010001010100" => A <= "000000000000000100"; -- Line 70   Column 5   Coefficient 0.00001526
         when "010001010101" => A <= "000000000000000000"; -- Line 70   Column 6   Coefficient 0.00000000
         when "010001010110" => A <= "000000000000000000"; -- Line 70   Column 7   Coefficient 0.00000000
         when "010001010111" => A <= "000000000000000000"; -- Line 70   Column 8   Coefficient 0.00000000
         when "010001011000" => A <= "000000000000000000"; -- Line 70   Column 9   Coefficient 0.00000000
         when "010001011001" => A <= "000000000000000000"; -- Line 70   Column 10   Coefficient 0.00000000
         when "010001011010" => A <= "000000000000000000"; -- Line 70   Column 11   Coefficient 0.00000000
         when "010001011011" => A <= "000000000000000000"; -- Line 70   Column 12   Coefficient 0.00000000
         when "010001011100" => A <= "000000000000000000"; -- Line 70   Column 13   Coefficient 0.00000000
         when "010001011101" => A <= "000000000000000000"; -- Line 70   Column 14   Coefficient 0.00000000
         when "010001011110" => A <= "111111111110010010"; -- Line 70   Column 15   Coefficient -0.00041962
         when "010001011111" => A <= "111110010000110000"; -- Line 70   Column 16   Coefficient -0.02716064
         when "010001100000" => A <= "001001000110101001"; -- Line 71   Column 1   Coefficient 0.14224625
         when "010001100001" => A <= "001000110101000000"; -- Line 71   Column 2   Coefficient 0.13793945
         when "010001100010" => A <= "111111100111100010"; -- Line 71   Column 3   Coefficient -0.00597382
         when "010001100011" => A <= "000000000010010011"; -- Line 71   Column 4   Coefficient 0.00056076
         when "010001100100" => A <= "000000000000000011"; -- Line 71   Column 5   Coefficient 0.00001144
         when "010001100101" => A <= "000000000000000000"; -- Line 71   Column 6   Coefficient 0.00000000
         when "010001100110" => A <= "000000000000000000"; -- Line 71   Column 7   Coefficient 0.00000000
         when "010001100111" => A <= "000000000000000000"; -- Line 71   Column 8   Coefficient 0.00000000
         when "010001101000" => A <= "000000000000000000"; -- Line 71   Column 9   Coefficient 0.00000000
         when "010001101001" => A <= "000000000000000000"; -- Line 71   Column 10   Coefficient 0.00000000
         when "010001101010" => A <= "000000000000000000"; -- Line 71   Column 11   Coefficient 0.00000000
         when "010001101011" => A <= "000000000000000000"; -- Line 71   Column 12   Coefficient 0.00000000
         when "010001101100" => A <= "000000000000000000"; -- Line 71   Column 13   Coefficient 0.00000000
         when "010001101101" => A <= "000000000000000000"; -- Line 71   Column 14   Coefficient 0.00000000
         when "010001101110" => A <= "111111111110100110"; -- Line 71   Column 15   Coefficient -0.00034332
         when "010001101111" => A <= "111110011011111010"; -- Line 71   Column 16   Coefficient -0.02443695
         when "010001110000" => A <= "000111100110110001"; -- Line 72   Column 1   Coefficient 0.11883926
         when "010001110001" => A <= "001010011001111000"; -- Line 72   Column 2   Coefficient 0.16256714
         when "010001110010" => A <= "111111010000101110"; -- Line 72   Column 3   Coefficient -0.01154327
         when "010001110011" => A <= "000000001001011000"; -- Line 72   Column 4   Coefficient 0.00228882
         when "010001110100" => A <= "111111111111110100"; -- Line 72   Column 5   Coefficient -0.00004578
         when "010001110101" => A <= "000000000000000000"; -- Line 72   Column 6   Coefficient 0.00000000
         when "010001110110" => A <= "000000000000000000"; -- Line 72   Column 7   Coefficient 0.00000000
         when "010001110111" => A <= "000000000000000000"; -- Line 72   Column 8   Coefficient 0.00000000
         when "010001111000" => A <= "000000000000000000"; -- Line 72   Column 9   Coefficient 0.00000000
         when "010001111001" => A <= "000000000000000000"; -- Line 72   Column 10   Coefficient 0.00000000
         when "010001111010" => A <= "000000000000000000"; -- Line 72   Column 11   Coefficient 0.00000000
         when "010001111011" => A <= "000000000000000000"; -- Line 72   Column 12   Coefficient 0.00000000
         when "010001111100" => A <= "000000000000000000"; -- Line 72   Column 13   Coefficient 0.00000000
         when "010001111101" => A <= "000000000000000000"; -- Line 72   Column 14   Coefficient 0.00000000
         when "010001111110" => A <= "111111111111001011"; -- Line 72   Column 15   Coefficient -0.00020218
         when "010001111111" => A <= "111110100110010011"; -- Line 72   Column 16   Coefficient -0.02190018
         when "010010000000" => A <= "000110000101110011"; -- Line 73   Column 1   Coefficient 0.09516525
         when "010010000001" => A <= "001011111101111010"; -- Line 73   Column 2   Coefficient 0.18698883
         when "010010000010" => A <= "111110111010000001"; -- Line 73   Column 3   Coefficient -0.01708603
         when "010010000011" => A <= "000000010001001000"; -- Line 73   Column 4   Coefficient 0.00418091
         when "010010000100" => A <= "111111111111100110"; -- Line 73   Column 5   Coefficient -0.00009918
         when "010010000101" => A <= "000000000000000000"; -- Line 73   Column 6   Coefficient 0.00000000
         when "010010000110" => A <= "000000000000000000"; -- Line 73   Column 7   Coefficient 0.00000000
         when "010010000111" => A <= "000000000000000000"; -- Line 73   Column 8   Coefficient 0.00000000
         when "010010001000" => A <= "000000000000000000"; -- Line 73   Column 9   Coefficient 0.00000000
         when "010010001001" => A <= "000000000000000000"; -- Line 73   Column 10   Coefficient 0.00000000
         when "010010001010" => A <= "000000000000000000"; -- Line 73   Column 11   Coefficient 0.00000000
         when "010010001011" => A <= "000000000000000000"; -- Line 73   Column 12   Coefficient 0.00000000
         when "010010001100" => A <= "000000000000000000"; -- Line 73   Column 13   Coefficient 0.00000000
         when "010010001101" => A <= "000000000000000000"; -- Line 73   Column 14   Coefficient 0.00000000
         when "010010001110" => A <= "000000000000000011"; -- Line 73   Column 15   Coefficient 0.00001144
         when "010010001111" => A <= "111110110001100001"; -- Line 73   Column 16   Coefficient -0.01916122
         when "010010010000" => A <= "000100010010000101"; -- Line 74   Column 1   Coefficient 0.06691360
         when "010010010001" => A <= "001101110100101001"; -- Line 74   Column 2   Coefficient 0.21597672
         when "010010010010" => A <= "111110011010010101"; -- Line 74   Column 3   Coefficient -0.02482224
         when "010010010011" => A <= "000000011001110100"; -- Line 74   Column 4   Coefficient 0.00630188
         when "010010010100" => A <= "000000000000000111"; -- Line 74   Column 5   Coefficient 0.00002670
         when "010010010101" => A <= "000000000000000000"; -- Line 74   Column 6   Coefficient 0.00000000
         when "010010010110" => A <= "000000000000000000"; -- Line 74   Column 7   Coefficient 0.00000000
         when "010010010111" => A <= "000000000000000000"; -- Line 74   Column 8   Coefficient 0.00000000
         when "010010011000" => A <= "000000000000000000"; -- Line 74   Column 9   Coefficient 0.00000000
         when "010010011001" => A <= "000000000000000000"; -- Line 74   Column 10   Coefficient 0.00000000
         when "010010011010" => A <= "000000000000000000"; -- Line 74   Column 11   Coefficient 0.00000000
         when "010010011011" => A <= "000000000000000000"; -- Line 74   Column 12   Coefficient 0.00000000
         when "010010011100" => A <= "000000000000000000"; -- Line 74   Column 13   Coefficient 0.00000000
         when "010010011101" => A <= "000000000000000000"; -- Line 74   Column 14   Coefficient 0.00000000
         when "010010011110" => A <= "000000000000001001"; -- Line 74   Column 15   Coefficient 0.00003433
         when "010010011111" => A <= "111111000100111001"; -- Line 74   Column 16   Coefficient -0.01443100
         when "010010100000" => A <= "000010011110111100"; -- Line 75   Column 1   Coefficient 0.03880310
         when "010010100001" => A <= "001111100101110011"; -- Line 75   Column 2   Coefficient 0.24360275
         when "010010100010" => A <= "111101111110110001"; -- Line 75   Column 3   Coefficient -0.03155136
         when "010010100011" => A <= "000000100001110011"; -- Line 75   Column 4   Coefficient 0.00825119
         when "010010100100" => A <= "000000000000110011"; -- Line 75   Column 5   Coefficient 0.00019455
         when "010010100101" => A <= "000000000000000000"; -- Line 75   Column 6   Coefficient 0.00000000
         when "010010100110" => A <= "000000000000000000"; -- Line 75   Column 7   Coefficient 0.00000000
         when "010010100111" => A <= "000000000000000000"; -- Line 75   Column 8   Coefficient 0.00000000
         when "010010101000" => A <= "000000000000000000"; -- Line 75   Column 9   Coefficient 0.00000000
         when "010010101001" => A <= "000000000000000000"; -- Line 75   Column 10   Coefficient 0.00000000
         when "010010101010" => A <= "000000000000000000"; -- Line 75   Column 11   Coefficient 0.00000000
         when "010010101011" => A <= "000000000000000000"; -- Line 75   Column 12   Coefficient 0.00000000
         when "010010101100" => A <= "000000000000000000"; -- Line 75   Column 13   Coefficient 0.00000000
         when "010010101101" => A <= "000000000000000000"; -- Line 75   Column 14   Coefficient 0.00000000
         when "010010101110" => A <= "000000000000000000"; -- Line 75   Column 15   Coefficient 0.00000000
         when "010010101111" => A <= "111111011001111001"; -- Line 75   Column 16   Coefficient -0.00930405
         when "010010110000" => A <= "000000100101011001"; -- Line 76   Column 1   Coefficient 0.00912857
         when "010010110001" => A <= "010001011110001011"; -- Line 76   Column 2   Coefficient 0.27299118
         when "010010110010" => A <= "111101011101101101"; -- Line 76   Column 3   Coefficient -0.03962326
         when "010010110011" => A <= "000000101011110101"; -- Line 76   Column 4   Coefficient 0.01070023
         when "010010110100" => A <= "000000000001100101"; -- Line 76   Column 5   Coefficient 0.00038528
         when "010010110101" => A <= "000000000000000000"; -- Line 76   Column 6   Coefficient 0.00000000
         when "010010110110" => A <= "000000000000000000"; -- Line 76   Column 7   Coefficient 0.00000000
         when "010010110111" => A <= "000000000000000000"; -- Line 76   Column 8   Coefficient 0.00000000
         when "010010111000" => A <= "000000000000000000"; -- Line 76   Column 9   Coefficient 0.00000000
         when "010010111001" => A <= "000000000000000000"; -- Line 76   Column 10   Coefficient 0.00000000
         when "010010111010" => A <= "000000000000000000"; -- Line 76   Column 11   Coefficient 0.00000000
         when "010010111011" => A <= "000000000000000000"; -- Line 76   Column 12   Coefficient 0.00000000
         when "010010111100" => A <= "000000000000000000"; -- Line 76   Column 13   Coefficient 0.00000000
         when "010010111101" => A <= "000000000000000000"; -- Line 76   Column 14   Coefficient 0.00000000
         when "010010111110" => A <= "000000000000000000"; -- Line 76   Column 15   Coefficient 0.00000000
         when "010010111111" => A <= "111111110001010101"; -- Line 76   Column 16   Coefficient -0.00358200
         when "010011000000" => A <= "111110110101100100"; -- Line 77   Column 1   Coefficient -0.01817322
         when "010011000001" => A <= "010011000101100111"; -- Line 77   Column 2   Coefficient 0.29824448
         when "010011000010" => A <= "111101000110110001"; -- Line 77   Column 3   Coefficient -0.04522324
         when "010011000011" => A <= "000000110100010110"; -- Line 77   Column 4   Coefficient 0.01277924
         when "010011000100" => A <= "000000000010010101"; -- Line 77   Column 5   Coefficient 0.00056839
         when "010011000101" => A <= "000000000000000000"; -- Line 77   Column 6   Coefficient 0.00000000
         when "010011000110" => A <= "000000000000000000"; -- Line 77   Column 7   Coefficient 0.00000000
         when "010011000111" => A <= "000000000000000000"; -- Line 77   Column 8   Coefficient 0.00000000
         when "010011001000" => A <= "000000000000000000"; -- Line 77   Column 9   Coefficient 0.00000000
         when "010011001001" => A <= "000000000000000000"; -- Line 77   Column 10   Coefficient 0.00000000
         when "010011001010" => A <= "000000000000000000"; -- Line 77   Column 11   Coefficient 0.00000000
         when "010011001011" => A <= "000000000000000000"; -- Line 77   Column 12   Coefficient 0.00000000
         when "010011001100" => A <= "000000000000000000"; -- Line 77   Column 13   Coefficient 0.00000000
         when "010011001101" => A <= "000000000000000000"; -- Line 77   Column 14   Coefficient 0.00000000
         when "010011001110" => A <= "000000000000000000"; -- Line 77   Column 15   Coefficient 0.00000000
         when "010011001111" => A <= "000000000111011010"; -- Line 77   Column 16   Coefficient 0.00180817
         when "010011010000" => A <= "111110000010011110"; -- Line 78   Column 1   Coefficient -0.03064728
         when "010011010001" => A <= "010011010010100110"; -- Line 78   Column 2   Coefficient 0.30141449
         when "010011010010" => A <= "111101100111001110"; -- Line 78   Column 3   Coefficient -0.03730011
         when "010011010011" => A <= "000000110010101110"; -- Line 78   Column 4   Coefficient 0.01238251
         when "010011010100" => A <= "000000000001111110"; -- Line 78   Column 5   Coefficient 0.00048065
         when "010011010101" => A <= "000000000000000000"; -- Line 78   Column 6   Coefficient 0.00000000
         when "010011010110" => A <= "000000000000000000"; -- Line 78   Column 7   Coefficient 0.00000000
         when "010011010111" => A <= "000000000000000000"; -- Line 78   Column 8   Coefficient 0.00000000
         when "010011011000" => A <= "000000000000000000"; -- Line 78   Column 9   Coefficient 0.00000000
         when "010011011001" => A <= "000000000000000000"; -- Line 78   Column 10   Coefficient 0.00000000
         when "010011011010" => A <= "000000000000000000"; -- Line 78   Column 11   Coefficient 0.00000000
         when "010011011011" => A <= "000000000000000000"; -- Line 78   Column 12   Coefficient 0.00000000
         when "010011011100" => A <= "000000000000000000"; -- Line 78   Column 13   Coefficient 0.00000000
         when "010011011101" => A <= "000000000000000000"; -- Line 78   Column 14   Coefficient 0.00000000
         when "010011011110" => A <= "000000000000000000"; -- Line 78   Column 15   Coefficient 0.00000000
         when "010011011111" => A <= "000000001111000010"; -- Line 78   Column 16   Coefficient 0.00366974
         when "010011100000" => A <= "111101101011101110"; -- Line 79   Column 1   Coefficient -0.03620148
         when "010011100001" => A <= "010010110100110100"; -- Line 79   Column 2   Coefficient 0.29414368
         when "010011100010" => A <= "111110100000101100"; -- Line 79   Column 3   Coefficient -0.02326965
         when "010011100011" => A <= "000000101101010111"; -- Line 79   Column 4   Coefficient 0.01107407
         when "010011100100" => A <= "000000000001000010"; -- Line 79   Column 5   Coefficient 0.00025177
         when "010011100101" => A <= "000000000000000000"; -- Line 79   Column 6   Coefficient 0.00000000
         when "010011100110" => A <= "000000000000000000"; -- Line 79   Column 7   Coefficient 0.00000000
         when "010011100111" => A <= "000000000000000000"; -- Line 79   Column 8   Coefficient 0.00000000
         when "010011101000" => A <= "000000000000000000"; -- Line 79   Column 9   Coefficient 0.00000000
         when "010011101001" => A <= "000000000000000000"; -- Line 79   Column 10   Coefficient 0.00000000
         when "010011101010" => A <= "000000000000000000"; -- Line 79   Column 11   Coefficient 0.00000000
         when "010011101011" => A <= "000000000000000000"; -- Line 79   Column 12   Coefficient 0.00000000
         when "010011101100" => A <= "000000000000000000"; -- Line 79   Column 13   Coefficient 0.00000000
         when "010011101101" => A <= "000000000000000000"; -- Line 79   Column 14   Coefficient 0.00000000
         when "010011101110" => A <= "000000000000000000"; -- Line 79   Column 15   Coefficient 0.00000000
         when "010011101111" => A <= "000000010000011000"; -- Line 79   Column 16   Coefficient 0.00399780
         when "010011110000" => A <= "111101100000101101"; -- Line 80   Column 1   Coefficient -0.03889084
         when "010011110001" => A <= "010010000001100011"; -- Line 80   Column 2   Coefficient 0.28162766
         when "010011110010" => A <= "111111101010001000"; -- Line 80   Column 3   Coefficient -0.00534058
         when "010011110011" => A <= "000000100010100100"; -- Line 80   Column 4   Coefficient 0.00843811
         when "010011110100" => A <= "000000000001001000"; -- Line 80   Column 5   Coefficient 0.00027466
         when "010011110101" => A <= "000000000000000000"; -- Line 80   Column 6   Coefficient 0.00000000
         when "010011110110" => A <= "000000000000000000"; -- Line 80   Column 7   Coefficient 0.00000000
         when "010011110111" => A <= "000000000000000000"; -- Line 80   Column 8   Coefficient 0.00000000
         when "010011111000" => A <= "000000000000000000"; -- Line 80   Column 9   Coefficient 0.00000000
         when "010011111001" => A <= "000000000000000000"; -- Line 80   Column 10   Coefficient 0.00000000
         when "010011111010" => A <= "000000000000000000"; -- Line 80   Column 11   Coefficient 0.00000000
         when "010011111011" => A <= "000000000000000000"; -- Line 80   Column 12   Coefficient 0.00000000
         when "010011111100" => A <= "000000000000000000"; -- Line 80   Column 13   Coefficient 0.00000000
         when "010011111101" => A <= "000000000000000000"; -- Line 80   Column 14   Coefficient 0.00000000
         when "010011111110" => A <= "000000000000000000"; -- Line 80   Column 15   Coefficient 0.00000000
         when "010011111111" => A <= "000000001111111100"; -- Line 80   Column 16   Coefficient 0.00389099
         when "010100000000" => A <= "111101100010001110"; -- Line 81   Column 1   Coefficient -0.03852081
         when "010100000001" => A <= "010000111010100101"; -- Line 81   Column 2   Coefficient 0.26430130
         when "010100000010" => A <= "000000111110100110"; -- Line 81   Column 3   Coefficient 0.01528168
         when "010100000011" => A <= "000000010110010000"; -- Line 81   Column 4   Coefficient 0.00543213
         when "010100000100" => A <= "000000000001001011"; -- Line 81   Column 5   Coefficient 0.00028610
         when "010100000101" => A <= "000000000000000000"; -- Line 81   Column 6   Coefficient 0.00000000
         when "010100000110" => A <= "000000000000000000"; -- Line 81   Column 7   Coefficient 0.00000000
         when "010100000111" => A <= "000000000000000000"; -- Line 81   Column 8   Coefficient 0.00000000
         when "010100001000" => A <= "000000000000000000"; -- Line 81   Column 9   Coefficient 0.00000000
         when "010100001001" => A <= "000000000000000000"; -- Line 81   Column 10   Coefficient 0.00000000
         when "010100001010" => A <= "000000000000000000"; -- Line 81   Column 11   Coefficient 0.00000000
         when "010100001011" => A <= "000000000000000000"; -- Line 81   Column 12   Coefficient 0.00000000
         when "010100001100" => A <= "000000000000000000"; -- Line 81   Column 13   Coefficient 0.00000000
         when "010100001101" => A <= "000000000000000000"; -- Line 81   Column 14   Coefficient 0.00000000
         when "010100001110" => A <= "000000000000000000"; -- Line 81   Column 15   Coefficient 0.00000000
         when "010100001111" => A <= "000000001101001100"; -- Line 81   Column 16   Coefficient 0.00321960
         when "010100010000" => A <= "111101100010101111"; -- Line 82   Column 1   Coefficient -0.03839493
         when "010100010001" => A <= "001111111010100001"; -- Line 82   Column 2   Coefficient 0.24866104
         when "010100010010" => A <= "000010000100001011"; -- Line 82   Column 3   Coefficient 0.03226852
         when "010100010011" => A <= "000000010100110111"; -- Line 82   Column 4   Coefficient 0.00509262
         when "010100010100" => A <= "111111111110110111"; -- Line 82   Column 5   Coefficient -0.00027847
         when "010100010101" => A <= "000000000000000000"; -- Line 82   Column 6   Coefficient 0.00000000
         when "010100010110" => A <= "000000000000000000"; -- Line 82   Column 7   Coefficient 0.00000000
         when "010100010111" => A <= "000000000000000000"; -- Line 82   Column 8   Coefficient 0.00000000
         when "010100011000" => A <= "000000000000000000"; -- Line 82   Column 9   Coefficient 0.00000000
         when "010100011001" => A <= "000000000000000000"; -- Line 82   Column 10   Coefficient 0.00000000
         when "010100011010" => A <= "000000000000000000"; -- Line 82   Column 11   Coefficient 0.00000000
         when "010100011011" => A <= "000000000000000000"; -- Line 82   Column 12   Coefficient 0.00000000
         when "010100011100" => A <= "000000000000000000"; -- Line 82   Column 13   Coefficient 0.00000000
         when "010100011101" => A <= "000000000000000000"; -- Line 82   Column 14   Coefficient 0.00000000
         when "010100011110" => A <= "000000000000000000"; -- Line 82   Column 15   Coefficient 0.00000000
         when "010100011111" => A <= "000000001010110110"; -- Line 82   Column 16   Coefficient 0.00264740
         when "010100100000" => A <= "111101100110110000"; -- Line 83   Column 1   Coefficient -0.03741455
         when "010100100001" => A <= "001110110101010100"; -- Line 83   Column 2   Coefficient 0.23176575
         when "010100100010" => A <= "000011001010010011"; -- Line 83   Column 3   Coefficient 0.04938889
         when "010100100011" => A <= "000000010100111001"; -- Line 83   Column 4   Coefficient 0.00510025
         when "010100100100" => A <= "111111111100011110"; -- Line 83   Column 5   Coefficient -0.00086212
         when "010100100101" => A <= "111111111111111111"; -- Line 83   Column 6   Coefficient -0.00000381
         when "010100100110" => A <= "000000000000000000"; -- Line 83   Column 7   Coefficient 0.00000000
         when "010100100111" => A <= "000000000000000000"; -- Line 83   Column 8   Coefficient 0.00000000
         when "010100101000" => A <= "000000000000000000"; -- Line 83   Column 9   Coefficient 0.00000000
         when "010100101001" => A <= "000000000000000000"; -- Line 83   Column 10   Coefficient 0.00000000
         when "010100101010" => A <= "000000000000000000"; -- Line 83   Column 11   Coefficient 0.00000000
         when "010100101011" => A <= "000000000000000000"; -- Line 83   Column 12   Coefficient 0.00000000
         when "010100101100" => A <= "000000000000000000"; -- Line 83   Column 13   Coefficient 0.00000000
         when "010100101101" => A <= "000000000000000000"; -- Line 83   Column 14   Coefficient 0.00000000
         when "010100101110" => A <= "000000000000000000"; -- Line 83   Column 15   Coefficient 0.00000000
         when "010100101111" => A <= "000000001000010011"; -- Line 83   Column 16   Coefficient 0.00202560
         when "010100110000" => A <= "111101110100001010"; -- Line 84   Column 1   Coefficient -0.03414154
         when "010100110001" => A <= "001101100011111111"; -- Line 84   Column 2   Coefficient 0.21191025
         when "010100110010" => A <= "000100010011001101"; -- Line 84   Column 3   Coefficient 0.06718826
         when "010100110011" => A <= "000000010111101010"; -- Line 84   Column 4   Coefficient 0.00577545
         when "010100110100" => A <= "111111111001000110"; -- Line 84   Column 5   Coefficient -0.00168610
         when "010100110101" => A <= "000000000000000011"; -- Line 84   Column 6   Coefficient 0.00001144
         when "010100110110" => A <= "000000000000000000"; -- Line 84   Column 7   Coefficient 0.00000000
         when "010100110111" => A <= "000000000000000000"; -- Line 84   Column 8   Coefficient 0.00000000
         when "010100111000" => A <= "000000000000000000"; -- Line 84   Column 9   Coefficient 0.00000000
         when "010100111001" => A <= "000000000000000000"; -- Line 84   Column 10   Coefficient 0.00000000
         when "010100111010" => A <= "000000000000000000"; -- Line 84   Column 11   Coefficient 0.00000000
         when "010100111011" => A <= "000000000000000000"; -- Line 84   Column 12   Coefficient 0.00000000
         when "010100111100" => A <= "000000000000000000"; -- Line 84   Column 13   Coefficient 0.00000000
         when "010100111101" => A <= "000000000000000000"; -- Line 84   Column 14   Coefficient 0.00000000
         when "010100111110" => A <= "000000000000000000"; -- Line 84   Column 15   Coefficient 0.00000000
         when "010100111111" => A <= "000000000011111000"; -- Line 84   Column 16   Coefficient 0.00094604
         when "010101000000" => A <= "111110000101010011"; -- Line 85   Column 1   Coefficient -0.02995682
         when "010101000001" => A <= "001100001011101000"; -- Line 85   Column 2   Coefficient 0.19033813
         when "010101000010" => A <= "000101100000010101"; -- Line 85   Column 3   Coefficient 0.08601761
         when "010101000011" => A <= "000000011000110111"; -- Line 85   Column 4   Coefficient 0.00606918
         when "010101000100" => A <= "111111110110011111"; -- Line 85   Column 5   Coefficient -0.00232315
         when "010101000101" => A <= "000000000000000110"; -- Line 85   Column 6   Coefficient 0.00002289
         when "010101000110" => A <= "000000000000000000"; -- Line 85   Column 7   Coefficient 0.00000000
         when "010101000111" => A <= "000000000000000000"; -- Line 85   Column 8   Coefficient 0.00000000
         when "010101001000" => A <= "000000000000000000"; -- Line 85   Column 9   Coefficient 0.00000000
         when "010101001001" => A <= "000000000000000000"; -- Line 85   Column 10   Coefficient 0.00000000
         when "010101001010" => A <= "000000000000000000"; -- Line 85   Column 11   Coefficient 0.00000000
         when "010101001011" => A <= "000000000000000000"; -- Line 85   Column 12   Coefficient 0.00000000
         when "010101001100" => A <= "000000000000000000"; -- Line 85   Column 13   Coefficient 0.00000000
         when "010101001101" => A <= "000000000000000000"; -- Line 85   Column 14   Coefficient 0.00000000
         when "010101001110" => A <= "000000000000000000"; -- Line 85   Column 15   Coefficient 0.00000000
         when "010101001111" => A <= "111111111111010011"; -- Line 85   Column 16   Coefficient -0.00017166
         when "010101010000" => A <= "111110010000110000"; -- Line 86   Column 1   Coefficient -0.02716064
         when "010101010001" => A <= "001010101100000111"; -- Line 86   Column 2   Coefficient 0.16701889
         when "010101010010" => A <= "000111000101010101"; -- Line 86   Column 3   Coefficient 0.11067581
         when "010101010011" => A <= "000000000100100100"; -- Line 86   Column 4   Coefficient 0.00111389
         when "010101010100" => A <= "111111111010111001"; -- Line 86   Column 5   Coefficient -0.00124741
         when "010101010101" => A <= "000000000000000100"; -- Line 86   Column 6   Coefficient 0.00001526
         when "010101010110" => A <= "000000000000000000"; -- Line 86   Column 7   Coefficient 0.00000000
         when "010101010111" => A <= "000000000000000000"; -- Line 86   Column 8   Coefficient 0.00000000
         when "010101011000" => A <= "000000000000000000"; -- Line 86   Column 9   Coefficient 0.00000000
         when "010101011001" => A <= "000000000000000000"; -- Line 86   Column 10   Coefficient 0.00000000
         when "010101011010" => A <= "000000000000000000"; -- Line 86   Column 11   Coefficient 0.00000000
         when "010101011011" => A <= "000000000000000000"; -- Line 86   Column 12   Coefficient 0.00000000
         when "010101011100" => A <= "000000000000000000"; -- Line 86   Column 13   Coefficient 0.00000000
         when "010101011101" => A <= "000000000000000000"; -- Line 86   Column 14   Coefficient 0.00000000
         when "010101011110" => A <= "000000000000000000"; -- Line 86   Column 15   Coefficient 0.00000000
         when "010101011111" => A <= "111111111110010010"; -- Line 86   Column 16   Coefficient -0.00041962
         when "010101100000" => A <= "111110011011111010"; -- Line 87   Column 1   Coefficient -0.02443695
         when "010101100001" => A <= "001001000110101001"; -- Line 87   Column 2   Coefficient 0.14224625
         when "010101100010" => A <= "001000110101000000"; -- Line 87   Column 3   Coefficient 0.13793945
         when "010101100011" => A <= "111111100111100010"; -- Line 87   Column 4   Coefficient -0.00597382
         when "010101100100" => A <= "000000000010010011"; -- Line 87   Column 5   Coefficient 0.00056076
         when "010101100101" => A <= "000000000000000011"; -- Line 87   Column 6   Coefficient 0.00001144
         when "010101100110" => A <= "000000000000000000"; -- Line 87   Column 7   Coefficient 0.00000000
         when "010101100111" => A <= "000000000000000000"; -- Line 87   Column 8   Coefficient 0.00000000
         when "010101101000" => A <= "000000000000000000"; -- Line 87   Column 9   Coefficient 0.00000000
         when "010101101001" => A <= "000000000000000000"; -- Line 87   Column 10   Coefficient 0.00000000
         when "010101101010" => A <= "000000000000000000"; -- Line 87   Column 11   Coefficient 0.00000000
         when "010101101011" => A <= "000000000000000000"; -- Line 87   Column 12   Coefficient 0.00000000
         when "010101101100" => A <= "000000000000000000"; -- Line 87   Column 13   Coefficient 0.00000000
         when "010101101101" => A <= "000000000000000000"; -- Line 87   Column 14   Coefficient 0.00000000
         when "010101101110" => A <= "000000000000000000"; -- Line 87   Column 15   Coefficient 0.00000000
         when "010101101111" => A <= "111111111110100110"; -- Line 87   Column 16   Coefficient -0.00034332
         when "010101110000" => A <= "111110100110010011"; -- Line 88   Column 1   Coefficient -0.02190018
         when "010101110001" => A <= "000111100110110001"; -- Line 88   Column 2   Coefficient 0.11883926
         when "010101110010" => A <= "001010011001111000"; -- Line 88   Column 3   Coefficient 0.16256714
         when "010101110011" => A <= "111111010000101110"; -- Line 88   Column 4   Coefficient -0.01154327
         when "010101110100" => A <= "000000001001011000"; -- Line 88   Column 5   Coefficient 0.00228882
         when "010101110101" => A <= "111111111111110100"; -- Line 88   Column 6   Coefficient -0.00004578
         when "010101110110" => A <= "000000000000000000"; -- Line 88   Column 7   Coefficient 0.00000000
         when "010101110111" => A <= "000000000000000000"; -- Line 88   Column 8   Coefficient 0.00000000
         when "010101111000" => A <= "000000000000000000"; -- Line 88   Column 9   Coefficient 0.00000000
         when "010101111001" => A <= "000000000000000000"; -- Line 88   Column 10   Coefficient 0.00000000
         when "010101111010" => A <= "000000000000000000"; -- Line 88   Column 11   Coefficient 0.00000000
         when "010101111011" => A <= "000000000000000000"; -- Line 88   Column 12   Coefficient 0.00000000
         when "010101111100" => A <= "000000000000000000"; -- Line 88   Column 13   Coefficient 0.00000000
         when "010101111101" => A <= "000000000000000000"; -- Line 88   Column 14   Coefficient 0.00000000
         when "010101111110" => A <= "000000000000000000"; -- Line 88   Column 15   Coefficient 0.00000000
         when "010101111111" => A <= "111111111111001011"; -- Line 88   Column 16   Coefficient -0.00020218
         when "010110000000" => A <= "111110110001100001"; -- Line 89   Column 1   Coefficient -0.01916122
         when "010110000001" => A <= "000110000101110011"; -- Line 89   Column 2   Coefficient 0.09516525
         when "010110000010" => A <= "001011111101111010"; -- Line 89   Column 3   Coefficient 0.18698883
         when "010110000011" => A <= "111110111010000001"; -- Line 89   Column 4   Coefficient -0.01708603
         when "010110000100" => A <= "000000010001001000"; -- Line 89   Column 5   Coefficient 0.00418091
         when "010110000101" => A <= "111111111111100110"; -- Line 89   Column 6   Coefficient -0.00009918
         when "010110000110" => A <= "000000000000000000"; -- Line 89   Column 7   Coefficient 0.00000000
         when "010110000111" => A <= "000000000000000000"; -- Line 89   Column 8   Coefficient 0.00000000
         when "010110001000" => A <= "000000000000000000"; -- Line 89   Column 9   Coefficient 0.00000000
         when "010110001001" => A <= "000000000000000000"; -- Line 89   Column 10   Coefficient 0.00000000
         when "010110001010" => A <= "000000000000000000"; -- Line 89   Column 11   Coefficient 0.00000000
         when "010110001011" => A <= "000000000000000000"; -- Line 89   Column 12   Coefficient 0.00000000
         when "010110001100" => A <= "000000000000000000"; -- Line 89   Column 13   Coefficient 0.00000000
         when "010110001101" => A <= "000000000000000000"; -- Line 89   Column 14   Coefficient 0.00000000
         when "010110001110" => A <= "000000000000000000"; -- Line 89   Column 15   Coefficient 0.00000000
         when "010110001111" => A <= "000000000000000011"; -- Line 89   Column 16   Coefficient 0.00001144
         when "010110010000" => A <= "111111000100111001"; -- Line 90   Column 1   Coefficient -0.01443100
         when "010110010001" => A <= "000100010010000101"; -- Line 90   Column 2   Coefficient 0.06691360
         when "010110010010" => A <= "001101110100101001"; -- Line 90   Column 3   Coefficient 0.21597672
         when "010110010011" => A <= "111110011010010101"; -- Line 90   Column 4   Coefficient -0.02482224
         when "010110010100" => A <= "000000011001110100"; -- Line 90   Column 5   Coefficient 0.00630188
         when "010110010101" => A <= "000000000000000111"; -- Line 90   Column 6   Coefficient 0.00002670
         when "010110010110" => A <= "000000000000000000"; -- Line 90   Column 7   Coefficient 0.00000000
         when "010110010111" => A <= "000000000000000000"; -- Line 90   Column 8   Coefficient 0.00000000
         when "010110011000" => A <= "000000000000000000"; -- Line 90   Column 9   Coefficient 0.00000000
         when "010110011001" => A <= "000000000000000000"; -- Line 90   Column 10   Coefficient 0.00000000
         when "010110011010" => A <= "000000000000000000"; -- Line 90   Column 11   Coefficient 0.00000000
         when "010110011011" => A <= "000000000000000000"; -- Line 90   Column 12   Coefficient 0.00000000
         when "010110011100" => A <= "000000000000000000"; -- Line 90   Column 13   Coefficient 0.00000000
         when "010110011101" => A <= "000000000000000000"; -- Line 90   Column 14   Coefficient 0.00000000
         when "010110011110" => A <= "000000000000000000"; -- Line 90   Column 15   Coefficient 0.00000000
         when "010110011111" => A <= "000000000000001001"; -- Line 90   Column 16   Coefficient 0.00003433
         when "010110100000" => A <= "111111011001111001"; -- Line 91   Column 1   Coefficient -0.00930405
         when "010110100001" => A <= "000010011110111100"; -- Line 91   Column 2   Coefficient 0.03880310
         when "010110100010" => A <= "001111100101110011"; -- Line 91   Column 3   Coefficient 0.24360275
         when "010110100011" => A <= "111101111110110001"; -- Line 91   Column 4   Coefficient -0.03155136
         when "010110100100" => A <= "000000100001110011"; -- Line 91   Column 5   Coefficient 0.00825119
         when "010110100101" => A <= "000000000000110011"; -- Line 91   Column 6   Coefficient 0.00019455
         when "010110100110" => A <= "000000000000000000"; -- Line 91   Column 7   Coefficient 0.00000000
         when "010110100111" => A <= "000000000000000000"; -- Line 91   Column 8   Coefficient 0.00000000
         when "010110101000" => A <= "000000000000000000"; -- Line 91   Column 9   Coefficient 0.00000000
         when "010110101001" => A <= "000000000000000000"; -- Line 91   Column 10   Coefficient 0.00000000
         when "010110101010" => A <= "000000000000000000"; -- Line 91   Column 11   Coefficient 0.00000000
         when "010110101011" => A <= "000000000000000000"; -- Line 91   Column 12   Coefficient 0.00000000
         when "010110101100" => A <= "000000000000000000"; -- Line 91   Column 13   Coefficient 0.00000000
         when "010110101101" => A <= "000000000000000000"; -- Line 91   Column 14   Coefficient 0.00000000
         when "010110101110" => A <= "000000000000000000"; -- Line 91   Column 15   Coefficient 0.00000000
         when "010110101111" => A <= "000000000000000000"; -- Line 91   Column 16   Coefficient 0.00000000
         when "010110110000" => A <= "111111110001010101"; -- Line 92   Column 1   Coefficient -0.00358200
         when "010110110001" => A <= "000000100101011001"; -- Line 92   Column 2   Coefficient 0.00912857
         when "010110110010" => A <= "010001011110001011"; -- Line 92   Column 3   Coefficient 0.27299118
         when "010110110011" => A <= "111101011101101101"; -- Line 92   Column 4   Coefficient -0.03962326
         when "010110110100" => A <= "000000101011110101"; -- Line 92   Column 5   Coefficient 0.01070023
         when "010110110101" => A <= "000000000001100101"; -- Line 92   Column 6   Coefficient 0.00038528
         when "010110110110" => A <= "000000000000000000"; -- Line 92   Column 7   Coefficient 0.00000000
         when "010110110111" => A <= "000000000000000000"; -- Line 92   Column 8   Coefficient 0.00000000
         when "010110111000" => A <= "000000000000000000"; -- Line 92   Column 9   Coefficient 0.00000000
         when "010110111001" => A <= "000000000000000000"; -- Line 92   Column 10   Coefficient 0.00000000
         when "010110111010" => A <= "000000000000000000"; -- Line 92   Column 11   Coefficient 0.00000000
         when "010110111011" => A <= "000000000000000000"; -- Line 92   Column 12   Coefficient 0.00000000
         when "010110111100" => A <= "000000000000000000"; -- Line 92   Column 13   Coefficient 0.00000000
         when "010110111101" => A <= "000000000000000000"; -- Line 92   Column 14   Coefficient 0.00000000
         when "010110111110" => A <= "000000000000000000"; -- Line 92   Column 15   Coefficient 0.00000000
         when "010110111111" => A <= "000000000000000000"; -- Line 92   Column 16   Coefficient 0.00000000
         when "010111000000" => A <= "000000000111011010"; -- Line 93   Column 1   Coefficient 0.00180817
         when "010111000001" => A <= "111110110101100100"; -- Line 93   Column 2   Coefficient -0.01817322
         when "010111000010" => A <= "010011000101100111"; -- Line 93   Column 3   Coefficient 0.29824448
         when "010111000011" => A <= "111101000110110001"; -- Line 93   Column 4   Coefficient -0.04522324
         when "010111000100" => A <= "000000110100010110"; -- Line 93   Column 5   Coefficient 0.01277924
         when "010111000101" => A <= "000000000010010101"; -- Line 93   Column 6   Coefficient 0.00056839
         when "010111000110" => A <= "000000000000000000"; -- Line 93   Column 7   Coefficient 0.00000000
         when "010111000111" => A <= "000000000000000000"; -- Line 93   Column 8   Coefficient 0.00000000
         when "010111001000" => A <= "000000000000000000"; -- Line 93   Column 9   Coefficient 0.00000000
         when "010111001001" => A <= "000000000000000000"; -- Line 93   Column 10   Coefficient 0.00000000
         when "010111001010" => A <= "000000000000000000"; -- Line 93   Column 11   Coefficient 0.00000000
         when "010111001011" => A <= "000000000000000000"; -- Line 93   Column 12   Coefficient 0.00000000
         when "010111001100" => A <= "000000000000000000"; -- Line 93   Column 13   Coefficient 0.00000000
         when "010111001101" => A <= "000000000000000000"; -- Line 93   Column 14   Coefficient 0.00000000
         when "010111001110" => A <= "000000000000000000"; -- Line 93   Column 15   Coefficient 0.00000000
         when "010111001111" => A <= "000000000000000000"; -- Line 93   Column 16   Coefficient 0.00000000
         when "010111010000" => A <= "000000001111000010"; -- Line 94   Column 1   Coefficient 0.00366974
         when "010111010001" => A <= "111110000010011110"; -- Line 94   Column 2   Coefficient -0.03064728
         when "010111010010" => A <= "010011010010100110"; -- Line 94   Column 3   Coefficient 0.30141449
         when "010111010011" => A <= "111101100111001110"; -- Line 94   Column 4   Coefficient -0.03730011
         when "010111010100" => A <= "000000110010101110"; -- Line 94   Column 5   Coefficient 0.01238251
         when "010111010101" => A <= "000000000001111110"; -- Line 94   Column 6   Coefficient 0.00048065
         when "010111010110" => A <= "000000000000000000"; -- Line 94   Column 7   Coefficient 0.00000000
         when "010111010111" => A <= "000000000000000000"; -- Line 94   Column 8   Coefficient 0.00000000
         when "010111011000" => A <= "000000000000000000"; -- Line 94   Column 9   Coefficient 0.00000000
         when "010111011001" => A <= "000000000000000000"; -- Line 94   Column 10   Coefficient 0.00000000
         when "010111011010" => A <= "000000000000000000"; -- Line 94   Column 11   Coefficient 0.00000000
         when "010111011011" => A <= "000000000000000000"; -- Line 94   Column 12   Coefficient 0.00000000
         when "010111011100" => A <= "000000000000000000"; -- Line 94   Column 13   Coefficient 0.00000000
         when "010111011101" => A <= "000000000000000000"; -- Line 94   Column 14   Coefficient 0.00000000
         when "010111011110" => A <= "000000000000000000"; -- Line 94   Column 15   Coefficient 0.00000000
         when "010111011111" => A <= "000000000000000000"; -- Line 94   Column 16   Coefficient 0.00000000
         when "010111100000" => A <= "000000010000011000"; -- Line 95   Column 1   Coefficient 0.00399780
         when "010111100001" => A <= "111101101011101110"; -- Line 95   Column 2   Coefficient -0.03620148
         when "010111100010" => A <= "010010110100110100"; -- Line 95   Column 3   Coefficient 0.29414368
         when "010111100011" => A <= "111110100000101100"; -- Line 95   Column 4   Coefficient -0.02326965
         when "010111100100" => A <= "000000101101010111"; -- Line 95   Column 5   Coefficient 0.01107407
         when "010111100101" => A <= "000000000001000010"; -- Line 95   Column 6   Coefficient 0.00025177
         when "010111100110" => A <= "000000000000000000"; -- Line 95   Column 7   Coefficient 0.00000000
         when "010111100111" => A <= "000000000000000000"; -- Line 95   Column 8   Coefficient 0.00000000
         when "010111101000" => A <= "000000000000000000"; -- Line 95   Column 9   Coefficient 0.00000000
         when "010111101001" => A <= "000000000000000000"; -- Line 95   Column 10   Coefficient 0.00000000
         when "010111101010" => A <= "000000000000000000"; -- Line 95   Column 11   Coefficient 0.00000000
         when "010111101011" => A <= "000000000000000000"; -- Line 95   Column 12   Coefficient 0.00000000
         when "010111101100" => A <= "000000000000000000"; -- Line 95   Column 13   Coefficient 0.00000000
         when "010111101101" => A <= "000000000000000000"; -- Line 95   Column 14   Coefficient 0.00000000
         when "010111101110" => A <= "000000000000000000"; -- Line 95   Column 15   Coefficient 0.00000000
         when "010111101111" => A <= "000000000000000000"; -- Line 95   Column 16   Coefficient 0.00000000
         when "010111110000" => A <= "000000001111111100"; -- Line 96   Column 1   Coefficient 0.00389099
         when "010111110001" => A <= "111101100000101101"; -- Line 96   Column 2   Coefficient -0.03889084
         when "010111110010" => A <= "010010000001100011"; -- Line 96   Column 3   Coefficient 0.28162766
         when "010111110011" => A <= "111111101010001000"; -- Line 96   Column 4   Coefficient -0.00534058
         when "010111110100" => A <= "000000100010100100"; -- Line 96   Column 5   Coefficient 0.00843811
         when "010111110101" => A <= "000000000001001000"; -- Line 96   Column 6   Coefficient 0.00027466
         when "010111110110" => A <= "000000000000000000"; -- Line 96   Column 7   Coefficient 0.00000000
         when "010111110111" => A <= "000000000000000000"; -- Line 96   Column 8   Coefficient 0.00000000
         when "010111111000" => A <= "000000000000000000"; -- Line 96   Column 9   Coefficient 0.00000000
         when "010111111001" => A <= "000000000000000000"; -- Line 96   Column 10   Coefficient 0.00000000
         when "010111111010" => A <= "000000000000000000"; -- Line 96   Column 11   Coefficient 0.00000000
         when "010111111011" => A <= "000000000000000000"; -- Line 96   Column 12   Coefficient 0.00000000
         when "010111111100" => A <= "000000000000000000"; -- Line 96   Column 13   Coefficient 0.00000000
         when "010111111101" => A <= "000000000000000000"; -- Line 96   Column 14   Coefficient 0.00000000
         when "010111111110" => A <= "000000000000000000"; -- Line 96   Column 15   Coefficient 0.00000000
         when "010111111111" => A <= "000000000000000000"; -- Line 96   Column 16   Coefficient 0.00000000
         when "011000000000" => A <= "000000001101001100"; -- Line 97   Column 1   Coefficient 0.00321960
         when "011000000001" => A <= "111101100010001110"; -- Line 97   Column 2   Coefficient -0.03852081
         when "011000000010" => A <= "010000111010100101"; -- Line 97   Column 3   Coefficient 0.26430130
         when "011000000011" => A <= "000000111110100110"; -- Line 97   Column 4   Coefficient 0.01528168
         when "011000000100" => A <= "000000010110010000"; -- Line 97   Column 5   Coefficient 0.00543213
         when "011000000101" => A <= "000000000001001011"; -- Line 97   Column 6   Coefficient 0.00028610
         when "011000000110" => A <= "000000000000000000"; -- Line 97   Column 7   Coefficient 0.00000000
         when "011000000111" => A <= "000000000000000000"; -- Line 97   Column 8   Coefficient 0.00000000
         when "011000001000" => A <= "000000000000000000"; -- Line 97   Column 9   Coefficient 0.00000000
         when "011000001001" => A <= "000000000000000000"; -- Line 97   Column 10   Coefficient 0.00000000
         when "011000001010" => A <= "000000000000000000"; -- Line 97   Column 11   Coefficient 0.00000000
         when "011000001011" => A <= "000000000000000000"; -- Line 97   Column 12   Coefficient 0.00000000
         when "011000001100" => A <= "000000000000000000"; -- Line 97   Column 13   Coefficient 0.00000000
         when "011000001101" => A <= "000000000000000000"; -- Line 97   Column 14   Coefficient 0.00000000
         when "011000001110" => A <= "000000000000000000"; -- Line 97   Column 15   Coefficient 0.00000000
         when "011000001111" => A <= "000000000000000000"; -- Line 97   Column 16   Coefficient 0.00000000
         when "011000010000" => A <= "000000001010110110"; -- Line 98   Column 1   Coefficient 0.00264740
         when "011000010001" => A <= "111101100010101111"; -- Line 98   Column 2   Coefficient -0.03839493
         when "011000010010" => A <= "001111111010100001"; -- Line 98   Column 3   Coefficient 0.24866104
         when "011000010011" => A <= "000010000100001011"; -- Line 98   Column 4   Coefficient 0.03226852
         when "011000010100" => A <= "000000010100110111"; -- Line 98   Column 5   Coefficient 0.00509262
         when "011000010101" => A <= "111111111110110111"; -- Line 98   Column 6   Coefficient -0.00027847
         when "011000010110" => A <= "000000000000000000"; -- Line 98   Column 7   Coefficient 0.00000000
         when "011000010111" => A <= "000000000000000000"; -- Line 98   Column 8   Coefficient 0.00000000
         when "011000011000" => A <= "000000000000000000"; -- Line 98   Column 9   Coefficient 0.00000000
         when "011000011001" => A <= "000000000000000000"; -- Line 98   Column 10   Coefficient 0.00000000
         when "011000011010" => A <= "000000000000000000"; -- Line 98   Column 11   Coefficient 0.00000000
         when "011000011011" => A <= "000000000000000000"; -- Line 98   Column 12   Coefficient 0.00000000
         when "011000011100" => A <= "000000000000000000"; -- Line 98   Column 13   Coefficient 0.00000000
         when "011000011101" => A <= "000000000000000000"; -- Line 98   Column 14   Coefficient 0.00000000
         when "011000011110" => A <= "000000000000000000"; -- Line 98   Column 15   Coefficient 0.00000000
         when "011000011111" => A <= "000000000000000000"; -- Line 98   Column 16   Coefficient 0.00000000
         when "011000100000" => A <= "000000001000010011"; -- Line 99   Column 1   Coefficient 0.00202560
         when "011000100001" => A <= "111101100110110000"; -- Line 99   Column 2   Coefficient -0.03741455
         when "011000100010" => A <= "001110110101010100"; -- Line 99   Column 3   Coefficient 0.23176575
         when "011000100011" => A <= "000011001010010011"; -- Line 99   Column 4   Coefficient 0.04938889
         when "011000100100" => A <= "000000010100111001"; -- Line 99   Column 5   Coefficient 0.00510025
         when "011000100101" => A <= "111111111100011110"; -- Line 99   Column 6   Coefficient -0.00086212
         when "011000100110" => A <= "111111111111111111"; -- Line 99   Column 7   Coefficient -0.00000381
         when "011000100111" => A <= "000000000000000000"; -- Line 99   Column 8   Coefficient 0.00000000
         when "011000101000" => A <= "000000000000000000"; -- Line 99   Column 9   Coefficient 0.00000000
         when "011000101001" => A <= "000000000000000000"; -- Line 99   Column 10   Coefficient 0.00000000
         when "011000101010" => A <= "000000000000000000"; -- Line 99   Column 11   Coefficient 0.00000000
         when "011000101011" => A <= "000000000000000000"; -- Line 99   Column 12   Coefficient 0.00000000
         when "011000101100" => A <= "000000000000000000"; -- Line 99   Column 13   Coefficient 0.00000000
         when "011000101101" => A <= "000000000000000000"; -- Line 99   Column 14   Coefficient 0.00000000
         when "011000101110" => A <= "000000000000000000"; -- Line 99   Column 15   Coefficient 0.00000000
         when "011000101111" => A <= "000000000000000000"; -- Line 99   Column 16   Coefficient 0.00000000
         when "011000110000" => A <= "000000000011111000"; -- Line 100   Column 1   Coefficient 0.00094604
         when "011000110001" => A <= "111101110100001010"; -- Line 100   Column 2   Coefficient -0.03414154
         when "011000110010" => A <= "001101100011111111"; -- Line 100   Column 3   Coefficient 0.21191025
         when "011000110011" => A <= "000100010011001101"; -- Line 100   Column 4   Coefficient 0.06718826
         when "011000110100" => A <= "000000010111101010"; -- Line 100   Column 5   Coefficient 0.00577545
         when "011000110101" => A <= "111111111001000110"; -- Line 100   Column 6   Coefficient -0.00168610
         when "011000110110" => A <= "000000000000000011"; -- Line 100   Column 7   Coefficient 0.00001144
         when "011000110111" => A <= "000000000000000000"; -- Line 100   Column 8   Coefficient 0.00000000
         when "011000111000" => A <= "000000000000000000"; -- Line 100   Column 9   Coefficient 0.00000000
         when "011000111001" => A <= "000000000000000000"; -- Line 100   Column 10   Coefficient 0.00000000
         when "011000111010" => A <= "000000000000000000"; -- Line 100   Column 11   Coefficient 0.00000000
         when "011000111011" => A <= "000000000000000000"; -- Line 100   Column 12   Coefficient 0.00000000
         when "011000111100" => A <= "000000000000000000"; -- Line 100   Column 13   Coefficient 0.00000000
         when "011000111101" => A <= "000000000000000000"; -- Line 100   Column 14   Coefficient 0.00000000
         when "011000111110" => A <= "000000000000000000"; -- Line 100   Column 15   Coefficient 0.00000000
         when "011000111111" => A <= "000000000000000000"; -- Line 100   Column 16   Coefficient 0.00000000
         when "011001000000" => A <= "111111111111010011"; -- Line 101   Column 1   Coefficient -0.00017166
         when "011001000001" => A <= "111110000101010011"; -- Line 101   Column 2   Coefficient -0.02995682
         when "011001000010" => A <= "001100001011101000"; -- Line 101   Column 3   Coefficient 0.19033813
         when "011001000011" => A <= "000101100000010101"; -- Line 101   Column 4   Coefficient 0.08601761
         when "011001000100" => A <= "000000011000110111"; -- Line 101   Column 5   Coefficient 0.00606918
         when "011001000101" => A <= "111111110110011111"; -- Line 101   Column 6   Coefficient -0.00232315
         when "011001000110" => A <= "000000000000000110"; -- Line 101   Column 7   Coefficient 0.00002289
         when "011001000111" => A <= "000000000000000000"; -- Line 101   Column 8   Coefficient 0.00000000
         when "011001001000" => A <= "000000000000000000"; -- Line 101   Column 9   Coefficient 0.00000000
         when "011001001001" => A <= "000000000000000000"; -- Line 101   Column 10   Coefficient 0.00000000
         when "011001001010" => A <= "000000000000000000"; -- Line 101   Column 11   Coefficient 0.00000000
         when "011001001011" => A <= "000000000000000000"; -- Line 101   Column 12   Coefficient 0.00000000
         when "011001001100" => A <= "000000000000000000"; -- Line 101   Column 13   Coefficient 0.00000000
         when "011001001101" => A <= "000000000000000000"; -- Line 101   Column 14   Coefficient 0.00000000
         when "011001001110" => A <= "000000000000000000"; -- Line 101   Column 15   Coefficient 0.00000000
         when "011001001111" => A <= "000000000000000000"; -- Line 101   Column 16   Coefficient 0.00000000
         when "011001010000" => A <= "111111111110010010"; -- Line 102   Column 1   Coefficient -0.00041962
         when "011001010001" => A <= "111110010000110000"; -- Line 102   Column 2   Coefficient -0.02716064
         when "011001010010" => A <= "001010101100000111"; -- Line 102   Column 3   Coefficient 0.16701889
         when "011001010011" => A <= "000111000101010101"; -- Line 102   Column 4   Coefficient 0.11067581
         when "011001010100" => A <= "000000000100100100"; -- Line 102   Column 5   Coefficient 0.00111389
         when "011001010101" => A <= "111111111010111001"; -- Line 102   Column 6   Coefficient -0.00124741
         when "011001010110" => A <= "000000000000000100"; -- Line 102   Column 7   Coefficient 0.00001526
         when "011001010111" => A <= "000000000000000000"; -- Line 102   Column 8   Coefficient 0.00000000
         when "011001011000" => A <= "000000000000000000"; -- Line 102   Column 9   Coefficient 0.00000000
         when "011001011001" => A <= "000000000000000000"; -- Line 102   Column 10   Coefficient 0.00000000
         when "011001011010" => A <= "000000000000000000"; -- Line 102   Column 11   Coefficient 0.00000000
         when "011001011011" => A <= "000000000000000000"; -- Line 102   Column 12   Coefficient 0.00000000
         when "011001011100" => A <= "000000000000000000"; -- Line 102   Column 13   Coefficient 0.00000000
         when "011001011101" => A <= "000000000000000000"; -- Line 102   Column 14   Coefficient 0.00000000
         when "011001011110" => A <= "000000000000000000"; -- Line 102   Column 15   Coefficient 0.00000000
         when "011001011111" => A <= "000000000000000000"; -- Line 102   Column 16   Coefficient 0.00000000
         when "011001100000" => A <= "111111111110100110"; -- Line 103   Column 1   Coefficient -0.00034332
         when "011001100001" => A <= "111110011011111010"; -- Line 103   Column 2   Coefficient -0.02443695
         when "011001100010" => A <= "001001000110101001"; -- Line 103   Column 3   Coefficient 0.14224625
         when "011001100011" => A <= "001000110101000000"; -- Line 103   Column 4   Coefficient 0.13793945
         when "011001100100" => A <= "111111100111100010"; -- Line 103   Column 5   Coefficient -0.00597382
         when "011001100101" => A <= "000000000010010011"; -- Line 103   Column 6   Coefficient 0.00056076
         when "011001100110" => A <= "000000000000000011"; -- Line 103   Column 7   Coefficient 0.00001144
         when "011001100111" => A <= "000000000000000000"; -- Line 103   Column 8   Coefficient 0.00000000
         when "011001101000" => A <= "000000000000000000"; -- Line 103   Column 9   Coefficient 0.00000000
         when "011001101001" => A <= "000000000000000000"; -- Line 103   Column 10   Coefficient 0.00000000
         when "011001101010" => A <= "000000000000000000"; -- Line 103   Column 11   Coefficient 0.00000000
         when "011001101011" => A <= "000000000000000000"; -- Line 103   Column 12   Coefficient 0.00000000
         when "011001101100" => A <= "000000000000000000"; -- Line 103   Column 13   Coefficient 0.00000000
         when "011001101101" => A <= "000000000000000000"; -- Line 103   Column 14   Coefficient 0.00000000
         when "011001101110" => A <= "000000000000000000"; -- Line 103   Column 15   Coefficient 0.00000000
         when "011001101111" => A <= "000000000000000000"; -- Line 103   Column 16   Coefficient 0.00000000
         when "011001110000" => A <= "111111111111001011"; -- Line 104   Column 1   Coefficient -0.00020218
         when "011001110001" => A <= "111110100110010011"; -- Line 104   Column 2   Coefficient -0.02190018
         when "011001110010" => A <= "000111100110110001"; -- Line 104   Column 3   Coefficient 0.11883926
         when "011001110011" => A <= "001010011001111000"; -- Line 104   Column 4   Coefficient 0.16256714
         when "011001110100" => A <= "111111010000101110"; -- Line 104   Column 5   Coefficient -0.01154327
         when "011001110101" => A <= "000000001001011000"; -- Line 104   Column 6   Coefficient 0.00228882
         when "011001110110" => A <= "111111111111110100"; -- Line 104   Column 7   Coefficient -0.00004578
         when "011001110111" => A <= "000000000000000000"; -- Line 104   Column 8   Coefficient 0.00000000
         when "011001111000" => A <= "000000000000000000"; -- Line 104   Column 9   Coefficient 0.00000000
         when "011001111001" => A <= "000000000000000000"; -- Line 104   Column 10   Coefficient 0.00000000
         when "011001111010" => A <= "000000000000000000"; -- Line 104   Column 11   Coefficient 0.00000000
         when "011001111011" => A <= "000000000000000000"; -- Line 104   Column 12   Coefficient 0.00000000
         when "011001111100" => A <= "000000000000000000"; -- Line 104   Column 13   Coefficient 0.00000000
         when "011001111101" => A <= "000000000000000000"; -- Line 104   Column 14   Coefficient 0.00000000
         when "011001111110" => A <= "000000000000000000"; -- Line 104   Column 15   Coefficient 0.00000000
         when "011001111111" => A <= "000000000000000000"; -- Line 104   Column 16   Coefficient 0.00000000
         when "011010000000" => A <= "000000000000000011"; -- Line 105   Column 1   Coefficient 0.00001144
         when "011010000001" => A <= "111110110001100001"; -- Line 105   Column 2   Coefficient -0.01916122
         when "011010000010" => A <= "000110000101110011"; -- Line 105   Column 3   Coefficient 0.09516525
         when "011010000011" => A <= "001011111101111010"; -- Line 105   Column 4   Coefficient 0.18698883
         when "011010000100" => A <= "111110111010000001"; -- Line 105   Column 5   Coefficient -0.01708603
         when "011010000101" => A <= "000000010001001000"; -- Line 105   Column 6   Coefficient 0.00418091
         when "011010000110" => A <= "111111111111100110"; -- Line 105   Column 7   Coefficient -0.00009918
         when "011010000111" => A <= "000000000000000000"; -- Line 105   Column 8   Coefficient 0.00000000
         when "011010001000" => A <= "000000000000000000"; -- Line 105   Column 9   Coefficient 0.00000000
         when "011010001001" => A <= "000000000000000000"; -- Line 105   Column 10   Coefficient 0.00000000
         when "011010001010" => A <= "000000000000000000"; -- Line 105   Column 11   Coefficient 0.00000000
         when "011010001011" => A <= "000000000000000000"; -- Line 105   Column 12   Coefficient 0.00000000
         when "011010001100" => A <= "000000000000000000"; -- Line 105   Column 13   Coefficient 0.00000000
         when "011010001101" => A <= "000000000000000000"; -- Line 105   Column 14   Coefficient 0.00000000
         when "011010001110" => A <= "000000000000000000"; -- Line 105   Column 15   Coefficient 0.00000000
         when "011010001111" => A <= "000000000000000000"; -- Line 105   Column 16   Coefficient 0.00000000
         when "011010010000" => A <= "000000000000001001"; -- Line 106   Column 1   Coefficient 0.00003433
         when "011010010001" => A <= "111111000100111001"; -- Line 106   Column 2   Coefficient -0.01443100
         when "011010010010" => A <= "000100010010000101"; -- Line 106   Column 3   Coefficient 0.06691360
         when "011010010011" => A <= "001101110100101001"; -- Line 106   Column 4   Coefficient 0.21597672
         when "011010010100" => A <= "111110011010010101"; -- Line 106   Column 5   Coefficient -0.02482224
         when "011010010101" => A <= "000000011001110100"; -- Line 106   Column 6   Coefficient 0.00630188
         when "011010010110" => A <= "000000000000000111"; -- Line 106   Column 7   Coefficient 0.00002670
         when "011010010111" => A <= "000000000000000000"; -- Line 106   Column 8   Coefficient 0.00000000
         when "011010011000" => A <= "000000000000000000"; -- Line 106   Column 9   Coefficient 0.00000000
         when "011010011001" => A <= "000000000000000000"; -- Line 106   Column 10   Coefficient 0.00000000
         when "011010011010" => A <= "000000000000000000"; -- Line 106   Column 11   Coefficient 0.00000000
         when "011010011011" => A <= "000000000000000000"; -- Line 106   Column 12   Coefficient 0.00000000
         when "011010011100" => A <= "000000000000000000"; -- Line 106   Column 13   Coefficient 0.00000000
         when "011010011101" => A <= "000000000000000000"; -- Line 106   Column 14   Coefficient 0.00000000
         when "011010011110" => A <= "000000000000000000"; -- Line 106   Column 15   Coefficient 0.00000000
         when "011010011111" => A <= "000000000000000000"; -- Line 106   Column 16   Coefficient 0.00000000
         when "011010100000" => A <= "000000000000000000"; -- Line 107   Column 1   Coefficient 0.00000000
         when "011010100001" => A <= "111111011001111001"; -- Line 107   Column 2   Coefficient -0.00930405
         when "011010100010" => A <= "000010011110111100"; -- Line 107   Column 3   Coefficient 0.03880310
         when "011010100011" => A <= "001111100101110011"; -- Line 107   Column 4   Coefficient 0.24360275
         when "011010100100" => A <= "111101111110110001"; -- Line 107   Column 5   Coefficient -0.03155136
         when "011010100101" => A <= "000000100001110011"; -- Line 107   Column 6   Coefficient 0.00825119
         when "011010100110" => A <= "000000000000110011"; -- Line 107   Column 7   Coefficient 0.00019455
         when "011010100111" => A <= "000000000000000000"; -- Line 107   Column 8   Coefficient 0.00000000
         when "011010101000" => A <= "000000000000000000"; -- Line 107   Column 9   Coefficient 0.00000000
         when "011010101001" => A <= "000000000000000000"; -- Line 107   Column 10   Coefficient 0.00000000
         when "011010101010" => A <= "000000000000000000"; -- Line 107   Column 11   Coefficient 0.00000000
         when "011010101011" => A <= "000000000000000000"; -- Line 107   Column 12   Coefficient 0.00000000
         when "011010101100" => A <= "000000000000000000"; -- Line 107   Column 13   Coefficient 0.00000000
         when "011010101101" => A <= "000000000000000000"; -- Line 107   Column 14   Coefficient 0.00000000
         when "011010101110" => A <= "000000000000000000"; -- Line 107   Column 15   Coefficient 0.00000000
         when "011010101111" => A <= "000000000000000000"; -- Line 107   Column 16   Coefficient 0.00000000
         when "011010110000" => A <= "000000000000000000"; -- Line 108   Column 1   Coefficient 0.00000000
         when "011010110001" => A <= "111111110001010101"; -- Line 108   Column 2   Coefficient -0.00358200
         when "011010110010" => A <= "000000100101011001"; -- Line 108   Column 3   Coefficient 0.00912857
         when "011010110011" => A <= "010001011110001011"; -- Line 108   Column 4   Coefficient 0.27299118
         when "011010110100" => A <= "111101011101101101"; -- Line 108   Column 5   Coefficient -0.03962326
         when "011010110101" => A <= "000000101011110101"; -- Line 108   Column 6   Coefficient 0.01070023
         when "011010110110" => A <= "000000000001100101"; -- Line 108   Column 7   Coefficient 0.00038528
         when "011010110111" => A <= "000000000000000000"; -- Line 108   Column 8   Coefficient 0.00000000
         when "011010111000" => A <= "000000000000000000"; -- Line 108   Column 9   Coefficient 0.00000000
         when "011010111001" => A <= "000000000000000000"; -- Line 108   Column 10   Coefficient 0.00000000
         when "011010111010" => A <= "000000000000000000"; -- Line 108   Column 11   Coefficient 0.00000000
         when "011010111011" => A <= "000000000000000000"; -- Line 108   Column 12   Coefficient 0.00000000
         when "011010111100" => A <= "000000000000000000"; -- Line 108   Column 13   Coefficient 0.00000000
         when "011010111101" => A <= "000000000000000000"; -- Line 108   Column 14   Coefficient 0.00000000
         when "011010111110" => A <= "000000000000000000"; -- Line 108   Column 15   Coefficient 0.00000000
         when "011010111111" => A <= "000000000000000000"; -- Line 108   Column 16   Coefficient 0.00000000
         when "011011000000" => A <= "000000000000000000"; -- Line 109   Column 1   Coefficient 0.00000000
         when "011011000001" => A <= "000000000111011010"; -- Line 109   Column 2   Coefficient 0.00180817
         when "011011000010" => A <= "111110110101100100"; -- Line 109   Column 3   Coefficient -0.01817322
         when "011011000011" => A <= "010011000101100111"; -- Line 109   Column 4   Coefficient 0.29824448
         when "011011000100" => A <= "111101000110110001"; -- Line 109   Column 5   Coefficient -0.04522324
         when "011011000101" => A <= "000000110100010110"; -- Line 109   Column 6   Coefficient 0.01277924
         when "011011000110" => A <= "000000000010010101"; -- Line 109   Column 7   Coefficient 0.00056839
         when "011011000111" => A <= "000000000000000000"; -- Line 109   Column 8   Coefficient 0.00000000
         when "011011001000" => A <= "000000000000000000"; -- Line 109   Column 9   Coefficient 0.00000000
         when "011011001001" => A <= "000000000000000000"; -- Line 109   Column 10   Coefficient 0.00000000
         when "011011001010" => A <= "000000000000000000"; -- Line 109   Column 11   Coefficient 0.00000000
         when "011011001011" => A <= "000000000000000000"; -- Line 109   Column 12   Coefficient 0.00000000
         when "011011001100" => A <= "000000000000000000"; -- Line 109   Column 13   Coefficient 0.00000000
         when "011011001101" => A <= "000000000000000000"; -- Line 109   Column 14   Coefficient 0.00000000
         when "011011001110" => A <= "000000000000000000"; -- Line 109   Column 15   Coefficient 0.00000000
         when "011011001111" => A <= "000000000000000000"; -- Line 109   Column 16   Coefficient 0.00000000
         when "011011010000" => A <= "000000000000000000"; -- Line 110   Column 1   Coefficient 0.00000000
         when "011011010001" => A <= "000000001111000010"; -- Line 110   Column 2   Coefficient 0.00366974
         when "011011010010" => A <= "111110000010011110"; -- Line 110   Column 3   Coefficient -0.03064728
         when "011011010011" => A <= "010011010010100110"; -- Line 110   Column 4   Coefficient 0.30141449
         when "011011010100" => A <= "111101100111001110"; -- Line 110   Column 5   Coefficient -0.03730011
         when "011011010101" => A <= "000000110010101110"; -- Line 110   Column 6   Coefficient 0.01238251
         when "011011010110" => A <= "000000000001111110"; -- Line 110   Column 7   Coefficient 0.00048065
         when "011011010111" => A <= "000000000000000000"; -- Line 110   Column 8   Coefficient 0.00000000
         when "011011011000" => A <= "000000000000000000"; -- Line 110   Column 9   Coefficient 0.00000000
         when "011011011001" => A <= "000000000000000000"; -- Line 110   Column 10   Coefficient 0.00000000
         when "011011011010" => A <= "000000000000000000"; -- Line 110   Column 11   Coefficient 0.00000000
         when "011011011011" => A <= "000000000000000000"; -- Line 110   Column 12   Coefficient 0.00000000
         when "011011011100" => A <= "000000000000000000"; -- Line 110   Column 13   Coefficient 0.00000000
         when "011011011101" => A <= "000000000000000000"; -- Line 110   Column 14   Coefficient 0.00000000
         when "011011011110" => A <= "000000000000000000"; -- Line 110   Column 15   Coefficient 0.00000000
         when "011011011111" => A <= "000000000000000000"; -- Line 110   Column 16   Coefficient 0.00000000
         when "011011100000" => A <= "000000000000000000"; -- Line 111   Column 1   Coefficient 0.00000000
         when "011011100001" => A <= "000000010000011000"; -- Line 111   Column 2   Coefficient 0.00399780
         when "011011100010" => A <= "111101101011101110"; -- Line 111   Column 3   Coefficient -0.03620148
         when "011011100011" => A <= "010010110100110100"; -- Line 111   Column 4   Coefficient 0.29414368
         when "011011100100" => A <= "111110100000101100"; -- Line 111   Column 5   Coefficient -0.02326965
         when "011011100101" => A <= "000000101101010111"; -- Line 111   Column 6   Coefficient 0.01107407
         when "011011100110" => A <= "000000000001000010"; -- Line 111   Column 7   Coefficient 0.00025177
         when "011011100111" => A <= "000000000000000000"; -- Line 111   Column 8   Coefficient 0.00000000
         when "011011101000" => A <= "000000000000000000"; -- Line 111   Column 9   Coefficient 0.00000000
         when "011011101001" => A <= "000000000000000000"; -- Line 111   Column 10   Coefficient 0.00000000
         when "011011101010" => A <= "000000000000000000"; -- Line 111   Column 11   Coefficient 0.00000000
         when "011011101011" => A <= "000000000000000000"; -- Line 111   Column 12   Coefficient 0.00000000
         when "011011101100" => A <= "000000000000000000"; -- Line 111   Column 13   Coefficient 0.00000000
         when "011011101101" => A <= "000000000000000000"; -- Line 111   Column 14   Coefficient 0.00000000
         when "011011101110" => A <= "000000000000000000"; -- Line 111   Column 15   Coefficient 0.00000000
         when "011011101111" => A <= "000000000000000000"; -- Line 111   Column 16   Coefficient 0.00000000
         when "011011110000" => A <= "000000000000000000"; -- Line 112   Column 1   Coefficient 0.00000000
         when "011011110001" => A <= "000000001111111100"; -- Line 112   Column 2   Coefficient 0.00389099
         when "011011110010" => A <= "111101100000101101"; -- Line 112   Column 3   Coefficient -0.03889084
         when "011011110011" => A <= "010010000001100011"; -- Line 112   Column 4   Coefficient 0.28162766
         when "011011110100" => A <= "111111101010001000"; -- Line 112   Column 5   Coefficient -0.00534058
         when "011011110101" => A <= "000000100010100100"; -- Line 112   Column 6   Coefficient 0.00843811
         when "011011110110" => A <= "000000000001001000"; -- Line 112   Column 7   Coefficient 0.00027466
         when "011011110111" => A <= "000000000000000000"; -- Line 112   Column 8   Coefficient 0.00000000
         when "011011111000" => A <= "000000000000000000"; -- Line 112   Column 9   Coefficient 0.00000000
         when "011011111001" => A <= "000000000000000000"; -- Line 112   Column 10   Coefficient 0.00000000
         when "011011111010" => A <= "000000000000000000"; -- Line 112   Column 11   Coefficient 0.00000000
         when "011011111011" => A <= "000000000000000000"; -- Line 112   Column 12   Coefficient 0.00000000
         when "011011111100" => A <= "000000000000000000"; -- Line 112   Column 13   Coefficient 0.00000000
         when "011011111101" => A <= "000000000000000000"; -- Line 112   Column 14   Coefficient 0.00000000
         when "011011111110" => A <= "000000000000000000"; -- Line 112   Column 15   Coefficient 0.00000000
         when "011011111111" => A <= "000000000000000000"; -- Line 112   Column 16   Coefficient 0.00000000
         when "011100000000" => A <= "000000000000000000"; -- Line 113   Column 1   Coefficient 0.00000000
         when "011100000001" => A <= "000000001101001100"; -- Line 113   Column 2   Coefficient 0.00321960
         when "011100000010" => A <= "111101100010001110"; -- Line 113   Column 3   Coefficient -0.03852081
         when "011100000011" => A <= "010000111010100101"; -- Line 113   Column 4   Coefficient 0.26430130
         when "011100000100" => A <= "000000111110100110"; -- Line 113   Column 5   Coefficient 0.01528168
         when "011100000101" => A <= "000000010110010000"; -- Line 113   Column 6   Coefficient 0.00543213
         when "011100000110" => A <= "000000000001001011"; -- Line 113   Column 7   Coefficient 0.00028610
         when "011100000111" => A <= "000000000000000000"; -- Line 113   Column 8   Coefficient 0.00000000
         when "011100001000" => A <= "000000000000000000"; -- Line 113   Column 9   Coefficient 0.00000000
         when "011100001001" => A <= "000000000000000000"; -- Line 113   Column 10   Coefficient 0.00000000
         when "011100001010" => A <= "000000000000000000"; -- Line 113   Column 11   Coefficient 0.00000000
         when "011100001011" => A <= "000000000000000000"; -- Line 113   Column 12   Coefficient 0.00000000
         when "011100001100" => A <= "000000000000000000"; -- Line 113   Column 13   Coefficient 0.00000000
         when "011100001101" => A <= "000000000000000000"; -- Line 113   Column 14   Coefficient 0.00000000
         when "011100001110" => A <= "000000000000000000"; -- Line 113   Column 15   Coefficient 0.00000000
         when "011100001111" => A <= "000000000000000000"; -- Line 113   Column 16   Coefficient 0.00000000
         when "011100010000" => A <= "000000000000000000"; -- Line 114   Column 1   Coefficient 0.00000000
         when "011100010001" => A <= "000000001010110110"; -- Line 114   Column 2   Coefficient 0.00264740
         when "011100010010" => A <= "111101100010101111"; -- Line 114   Column 3   Coefficient -0.03839493
         when "011100010011" => A <= "001111111010100001"; -- Line 114   Column 4   Coefficient 0.24866104
         when "011100010100" => A <= "000010000100001011"; -- Line 114   Column 5   Coefficient 0.03226852
         when "011100010101" => A <= "000000010100110111"; -- Line 114   Column 6   Coefficient 0.00509262
         when "011100010110" => A <= "111111111110110111"; -- Line 114   Column 7   Coefficient -0.00027847
         when "011100010111" => A <= "000000000000000000"; -- Line 114   Column 8   Coefficient 0.00000000
         when "011100011000" => A <= "000000000000000000"; -- Line 114   Column 9   Coefficient 0.00000000
         when "011100011001" => A <= "000000000000000000"; -- Line 114   Column 10   Coefficient 0.00000000
         when "011100011010" => A <= "000000000000000000"; -- Line 114   Column 11   Coefficient 0.00000000
         when "011100011011" => A <= "000000000000000000"; -- Line 114   Column 12   Coefficient 0.00000000
         when "011100011100" => A <= "000000000000000000"; -- Line 114   Column 13   Coefficient 0.00000000
         when "011100011101" => A <= "000000000000000000"; -- Line 114   Column 14   Coefficient 0.00000000
         when "011100011110" => A <= "000000000000000000"; -- Line 114   Column 15   Coefficient 0.00000000
         when "011100011111" => A <= "000000000000000000"; -- Line 114   Column 16   Coefficient 0.00000000
         when "011100100000" => A <= "000000000000000000"; -- Line 115   Column 1   Coefficient 0.00000000
         when "011100100001" => A <= "000000001000010011"; -- Line 115   Column 2   Coefficient 0.00202560
         when "011100100010" => A <= "111101100110110000"; -- Line 115   Column 3   Coefficient -0.03741455
         when "011100100011" => A <= "001110110101010100"; -- Line 115   Column 4   Coefficient 0.23176575
         when "011100100100" => A <= "000011001010010011"; -- Line 115   Column 5   Coefficient 0.04938889
         when "011100100101" => A <= "000000010100111001"; -- Line 115   Column 6   Coefficient 0.00510025
         when "011100100110" => A <= "111111111100011110"; -- Line 115   Column 7   Coefficient -0.00086212
         when "011100100111" => A <= "111111111111111111"; -- Line 115   Column 8   Coefficient -0.00000381
         when "011100101000" => A <= "000000000000000000"; -- Line 115   Column 9   Coefficient 0.00000000
         when "011100101001" => A <= "000000000000000000"; -- Line 115   Column 10   Coefficient 0.00000000
         when "011100101010" => A <= "000000000000000000"; -- Line 115   Column 11   Coefficient 0.00000000
         when "011100101011" => A <= "000000000000000000"; -- Line 115   Column 12   Coefficient 0.00000000
         when "011100101100" => A <= "000000000000000000"; -- Line 115   Column 13   Coefficient 0.00000000
         when "011100101101" => A <= "000000000000000000"; -- Line 115   Column 14   Coefficient 0.00000000
         when "011100101110" => A <= "000000000000000000"; -- Line 115   Column 15   Coefficient 0.00000000
         when "011100101111" => A <= "000000000000000000"; -- Line 115   Column 16   Coefficient 0.00000000
         when "011100110000" => A <= "000000000000000000"; -- Line 116   Column 1   Coefficient 0.00000000
         when "011100110001" => A <= "000000000011111000"; -- Line 116   Column 2   Coefficient 0.00094604
         when "011100110010" => A <= "111101110100001010"; -- Line 116   Column 3   Coefficient -0.03414154
         when "011100110011" => A <= "001101100011111111"; -- Line 116   Column 4   Coefficient 0.21191025
         when "011100110100" => A <= "000100010011001101"; -- Line 116   Column 5   Coefficient 0.06718826
         when "011100110101" => A <= "000000010111101010"; -- Line 116   Column 6   Coefficient 0.00577545
         when "011100110110" => A <= "111111111001000110"; -- Line 116   Column 7   Coefficient -0.00168610
         when "011100110111" => A <= "000000000000000011"; -- Line 116   Column 8   Coefficient 0.00001144
         when "011100111000" => A <= "000000000000000000"; -- Line 116   Column 9   Coefficient 0.00000000
         when "011100111001" => A <= "000000000000000000"; -- Line 116   Column 10   Coefficient 0.00000000
         when "011100111010" => A <= "000000000000000000"; -- Line 116   Column 11   Coefficient 0.00000000
         when "011100111011" => A <= "000000000000000000"; -- Line 116   Column 12   Coefficient 0.00000000
         when "011100111100" => A <= "000000000000000000"; -- Line 116   Column 13   Coefficient 0.00000000
         when "011100111101" => A <= "000000000000000000"; -- Line 116   Column 14   Coefficient 0.00000000
         when "011100111110" => A <= "000000000000000000"; -- Line 116   Column 15   Coefficient 0.00000000
         when "011100111111" => A <= "000000000000000000"; -- Line 116   Column 16   Coefficient 0.00000000
         when "011101000000" => A <= "000000000000000000"; -- Line 117   Column 1   Coefficient 0.00000000
         when "011101000001" => A <= "111111111111010011"; -- Line 117   Column 2   Coefficient -0.00017166
         when "011101000010" => A <= "111110000101010011"; -- Line 117   Column 3   Coefficient -0.02995682
         when "011101000011" => A <= "001100001011101000"; -- Line 117   Column 4   Coefficient 0.19033813
         when "011101000100" => A <= "000101100000010101"; -- Line 117   Column 5   Coefficient 0.08601761
         when "011101000101" => A <= "000000011000110111"; -- Line 117   Column 6   Coefficient 0.00606918
         when "011101000110" => A <= "111111110110011111"; -- Line 117   Column 7   Coefficient -0.00232315
         when "011101000111" => A <= "000000000000000110"; -- Line 117   Column 8   Coefficient 0.00002289
         when "011101001000" => A <= "000000000000000000"; -- Line 117   Column 9   Coefficient 0.00000000
         when "011101001001" => A <= "000000000000000000"; -- Line 117   Column 10   Coefficient 0.00000000
         when "011101001010" => A <= "000000000000000000"; -- Line 117   Column 11   Coefficient 0.00000000
         when "011101001011" => A <= "000000000000000000"; -- Line 117   Column 12   Coefficient 0.00000000
         when "011101001100" => A <= "000000000000000000"; -- Line 117   Column 13   Coefficient 0.00000000
         when "011101001101" => A <= "000000000000000000"; -- Line 117   Column 14   Coefficient 0.00000000
         when "011101001110" => A <= "000000000000000000"; -- Line 117   Column 15   Coefficient 0.00000000
         when "011101001111" => A <= "000000000000000000"; -- Line 117   Column 16   Coefficient 0.00000000
         when "011101010000" => A <= "000000000000000000"; -- Line 118   Column 1   Coefficient 0.00000000
         when "011101010001" => A <= "111111111110010010"; -- Line 118   Column 2   Coefficient -0.00041962
         when "011101010010" => A <= "111110010000110000"; -- Line 118   Column 3   Coefficient -0.02716064
         when "011101010011" => A <= "001010101100000111"; -- Line 118   Column 4   Coefficient 0.16701889
         when "011101010100" => A <= "000111000101010101"; -- Line 118   Column 5   Coefficient 0.11067581
         when "011101010101" => A <= "000000000100100100"; -- Line 118   Column 6   Coefficient 0.00111389
         when "011101010110" => A <= "111111111010111001"; -- Line 118   Column 7   Coefficient -0.00124741
         when "011101010111" => A <= "000000000000000100"; -- Line 118   Column 8   Coefficient 0.00001526
         when "011101011000" => A <= "000000000000000000"; -- Line 118   Column 9   Coefficient 0.00000000
         when "011101011001" => A <= "000000000000000000"; -- Line 118   Column 10   Coefficient 0.00000000
         when "011101011010" => A <= "000000000000000000"; -- Line 118   Column 11   Coefficient 0.00000000
         when "011101011011" => A <= "000000000000000000"; -- Line 118   Column 12   Coefficient 0.00000000
         when "011101011100" => A <= "000000000000000000"; -- Line 118   Column 13   Coefficient 0.00000000
         when "011101011101" => A <= "000000000000000000"; -- Line 118   Column 14   Coefficient 0.00000000
         when "011101011110" => A <= "000000000000000000"; -- Line 118   Column 15   Coefficient 0.00000000
         when "011101011111" => A <= "000000000000000000"; -- Line 118   Column 16   Coefficient 0.00000000
         when "011101100000" => A <= "000000000000000000"; -- Line 119   Column 1   Coefficient 0.00000000
         when "011101100001" => A <= "111111111110100110"; -- Line 119   Column 2   Coefficient -0.00034332
         when "011101100010" => A <= "111110011011111010"; -- Line 119   Column 3   Coefficient -0.02443695
         when "011101100011" => A <= "001001000110101001"; -- Line 119   Column 4   Coefficient 0.14224625
         when "011101100100" => A <= "001000110101000000"; -- Line 119   Column 5   Coefficient 0.13793945
         when "011101100101" => A <= "111111100111100010"; -- Line 119   Column 6   Coefficient -0.00597382
         when "011101100110" => A <= "000000000010010011"; -- Line 119   Column 7   Coefficient 0.00056076
         when "011101100111" => A <= "000000000000000011"; -- Line 119   Column 8   Coefficient 0.00001144
         when "011101101000" => A <= "000000000000000000"; -- Line 119   Column 9   Coefficient 0.00000000
         when "011101101001" => A <= "000000000000000000"; -- Line 119   Column 10   Coefficient 0.00000000
         when "011101101010" => A <= "000000000000000000"; -- Line 119   Column 11   Coefficient 0.00000000
         when "011101101011" => A <= "000000000000000000"; -- Line 119   Column 12   Coefficient 0.00000000
         when "011101101100" => A <= "000000000000000000"; -- Line 119   Column 13   Coefficient 0.00000000
         when "011101101101" => A <= "000000000000000000"; -- Line 119   Column 14   Coefficient 0.00000000
         when "011101101110" => A <= "000000000000000000"; -- Line 119   Column 15   Coefficient 0.00000000
         when "011101101111" => A <= "000000000000000000"; -- Line 119   Column 16   Coefficient 0.00000000
         when "011101110000" => A <= "000000000000000000"; -- Line 120   Column 1   Coefficient 0.00000000
         when "011101110001" => A <= "111111111111001011"; -- Line 120   Column 2   Coefficient -0.00020218
         when "011101110010" => A <= "111110100110010011"; -- Line 120   Column 3   Coefficient -0.02190018
         when "011101110011" => A <= "000111100110110001"; -- Line 120   Column 4   Coefficient 0.11883926
         when "011101110100" => A <= "001010011001111000"; -- Line 120   Column 5   Coefficient 0.16256714
         when "011101110101" => A <= "111111010000101110"; -- Line 120   Column 6   Coefficient -0.01154327
         when "011101110110" => A <= "000000001001011000"; -- Line 120   Column 7   Coefficient 0.00228882
         when "011101110111" => A <= "111111111111110100"; -- Line 120   Column 8   Coefficient -0.00004578
         when "011101111000" => A <= "000000000000000000"; -- Line 120   Column 9   Coefficient 0.00000000
         when "011101111001" => A <= "000000000000000000"; -- Line 120   Column 10   Coefficient 0.00000000
         when "011101111010" => A <= "000000000000000000"; -- Line 120   Column 11   Coefficient 0.00000000
         when "011101111011" => A <= "000000000000000000"; -- Line 120   Column 12   Coefficient 0.00000000
         when "011101111100" => A <= "000000000000000000"; -- Line 120   Column 13   Coefficient 0.00000000
         when "011101111101" => A <= "000000000000000000"; -- Line 120   Column 14   Coefficient 0.00000000
         when "011101111110" => A <= "000000000000000000"; -- Line 120   Column 15   Coefficient 0.00000000
         when "011101111111" => A <= "000000000000000000"; -- Line 120   Column 16   Coefficient 0.00000000
         when "011110000000" => A <= "000000000000000000"; -- Line 121   Column 1   Coefficient 0.00000000
         when "011110000001" => A <= "000000000000000011"; -- Line 121   Column 2   Coefficient 0.00001144
         when "011110000010" => A <= "111110110001100001"; -- Line 121   Column 3   Coefficient -0.01916122
         when "011110000011" => A <= "000110000101110011"; -- Line 121   Column 4   Coefficient 0.09516525
         when "011110000100" => A <= "001011111101111010"; -- Line 121   Column 5   Coefficient 0.18698883
         when "011110000101" => A <= "111110111010000001"; -- Line 121   Column 6   Coefficient -0.01708603
         when "011110000110" => A <= "000000010001001000"; -- Line 121   Column 7   Coefficient 0.00418091
         when "011110000111" => A <= "111111111111100110"; -- Line 121   Column 8   Coefficient -0.00009918
         when "011110001000" => A <= "000000000000000000"; -- Line 121   Column 9   Coefficient 0.00000000
         when "011110001001" => A <= "000000000000000000"; -- Line 121   Column 10   Coefficient 0.00000000
         when "011110001010" => A <= "000000000000000000"; -- Line 121   Column 11   Coefficient 0.00000000
         when "011110001011" => A <= "000000000000000000"; -- Line 121   Column 12   Coefficient 0.00000000
         when "011110001100" => A <= "000000000000000000"; -- Line 121   Column 13   Coefficient 0.00000000
         when "011110001101" => A <= "000000000000000000"; -- Line 121   Column 14   Coefficient 0.00000000
         when "011110001110" => A <= "000000000000000000"; -- Line 121   Column 15   Coefficient 0.00000000
         when "011110001111" => A <= "000000000000000000"; -- Line 121   Column 16   Coefficient 0.00000000
         when "011110010000" => A <= "000000000000000000"; -- Line 122   Column 1   Coefficient 0.00000000
         when "011110010001" => A <= "000000000000001001"; -- Line 122   Column 2   Coefficient 0.00003433
         when "011110010010" => A <= "111111000100111001"; -- Line 122   Column 3   Coefficient -0.01443100
         when "011110010011" => A <= "000100010010000101"; -- Line 122   Column 4   Coefficient 0.06691360
         when "011110010100" => A <= "001101110100101001"; -- Line 122   Column 5   Coefficient 0.21597672
         when "011110010101" => A <= "111110011010010101"; -- Line 122   Column 6   Coefficient -0.02482224
         when "011110010110" => A <= "000000011001110100"; -- Line 122   Column 7   Coefficient 0.00630188
         when "011110010111" => A <= "000000000000000111"; -- Line 122   Column 8   Coefficient 0.00002670
         when "011110011000" => A <= "000000000000000000"; -- Line 122   Column 9   Coefficient 0.00000000
         when "011110011001" => A <= "000000000000000000"; -- Line 122   Column 10   Coefficient 0.00000000
         when "011110011010" => A <= "000000000000000000"; -- Line 122   Column 11   Coefficient 0.00000000
         when "011110011011" => A <= "000000000000000000"; -- Line 122   Column 12   Coefficient 0.00000000
         when "011110011100" => A <= "000000000000000000"; -- Line 122   Column 13   Coefficient 0.00000000
         when "011110011101" => A <= "000000000000000000"; -- Line 122   Column 14   Coefficient 0.00000000
         when "011110011110" => A <= "000000000000000000"; -- Line 122   Column 15   Coefficient 0.00000000
         when "011110011111" => A <= "000000000000000000"; -- Line 122   Column 16   Coefficient 0.00000000
         when "011110100000" => A <= "000000000000000000"; -- Line 123   Column 1   Coefficient 0.00000000
         when "011110100001" => A <= "000000000000000000"; -- Line 123   Column 2   Coefficient 0.00000000
         when "011110100010" => A <= "111111011001111001"; -- Line 123   Column 3   Coefficient -0.00930405
         when "011110100011" => A <= "000010011110111100"; -- Line 123   Column 4   Coefficient 0.03880310
         when "011110100100" => A <= "001111100101110011"; -- Line 123   Column 5   Coefficient 0.24360275
         when "011110100101" => A <= "111101111110110001"; -- Line 123   Column 6   Coefficient -0.03155136
         when "011110100110" => A <= "000000100001110011"; -- Line 123   Column 7   Coefficient 0.00825119
         when "011110100111" => A <= "000000000000110011"; -- Line 123   Column 8   Coefficient 0.00019455
         when "011110101000" => A <= "000000000000000000"; -- Line 123   Column 9   Coefficient 0.00000000
         when "011110101001" => A <= "000000000000000000"; -- Line 123   Column 10   Coefficient 0.00000000
         when "011110101010" => A <= "000000000000000000"; -- Line 123   Column 11   Coefficient 0.00000000
         when "011110101011" => A <= "000000000000000000"; -- Line 123   Column 12   Coefficient 0.00000000
         when "011110101100" => A <= "000000000000000000"; -- Line 123   Column 13   Coefficient 0.00000000
         when "011110101101" => A <= "000000000000000000"; -- Line 123   Column 14   Coefficient 0.00000000
         when "011110101110" => A <= "000000000000000000"; -- Line 123   Column 15   Coefficient 0.00000000
         when "011110101111" => A <= "000000000000000000"; -- Line 123   Column 16   Coefficient 0.00000000
         when "011110110000" => A <= "000000000000000000"; -- Line 124   Column 1   Coefficient 0.00000000
         when "011110110001" => A <= "000000000000000000"; -- Line 124   Column 2   Coefficient 0.00000000
         when "011110110010" => A <= "111111110001010101"; -- Line 124   Column 3   Coefficient -0.00358200
         when "011110110011" => A <= "000000100101011001"; -- Line 124   Column 4   Coefficient 0.00912857
         when "011110110100" => A <= "010001011110001011"; -- Line 124   Column 5   Coefficient 0.27299118
         when "011110110101" => A <= "111101011101101101"; -- Line 124   Column 6   Coefficient -0.03962326
         when "011110110110" => A <= "000000101011110101"; -- Line 124   Column 7   Coefficient 0.01070023
         when "011110110111" => A <= "000000000001100101"; -- Line 124   Column 8   Coefficient 0.00038528
         when "011110111000" => A <= "000000000000000000"; -- Line 124   Column 9   Coefficient 0.00000000
         when "011110111001" => A <= "000000000000000000"; -- Line 124   Column 10   Coefficient 0.00000000
         when "011110111010" => A <= "000000000000000000"; -- Line 124   Column 11   Coefficient 0.00000000
         when "011110111011" => A <= "000000000000000000"; -- Line 124   Column 12   Coefficient 0.00000000
         when "011110111100" => A <= "000000000000000000"; -- Line 124   Column 13   Coefficient 0.00000000
         when "011110111101" => A <= "000000000000000000"; -- Line 124   Column 14   Coefficient 0.00000000
         when "011110111110" => A <= "000000000000000000"; -- Line 124   Column 15   Coefficient 0.00000000
         when "011110111111" => A <= "000000000000000000"; -- Line 124   Column 16   Coefficient 0.00000000
         when "011111000000" => A <= "000000000000000000"; -- Line 125   Column 1   Coefficient 0.00000000
         when "011111000001" => A <= "000000000000000000"; -- Line 125   Column 2   Coefficient 0.00000000
         when "011111000010" => A <= "000000000111011010"; -- Line 125   Column 3   Coefficient 0.00180817
         when "011111000011" => A <= "111110110101100100"; -- Line 125   Column 4   Coefficient -0.01817322
         when "011111000100" => A <= "010011000101100111"; -- Line 125   Column 5   Coefficient 0.29824448
         when "011111000101" => A <= "111101000110110001"; -- Line 125   Column 6   Coefficient -0.04522324
         when "011111000110" => A <= "000000110100010110"; -- Line 125   Column 7   Coefficient 0.01277924
         when "011111000111" => A <= "000000000010010101"; -- Line 125   Column 8   Coefficient 0.00056839
         when "011111001000" => A <= "000000000000000000"; -- Line 125   Column 9   Coefficient 0.00000000
         when "011111001001" => A <= "000000000000000000"; -- Line 125   Column 10   Coefficient 0.00000000
         when "011111001010" => A <= "000000000000000000"; -- Line 125   Column 11   Coefficient 0.00000000
         when "011111001011" => A <= "000000000000000000"; -- Line 125   Column 12   Coefficient 0.00000000
         when "011111001100" => A <= "000000000000000000"; -- Line 125   Column 13   Coefficient 0.00000000
         when "011111001101" => A <= "000000000000000000"; -- Line 125   Column 14   Coefficient 0.00000000
         when "011111001110" => A <= "000000000000000000"; -- Line 125   Column 15   Coefficient 0.00000000
         when "011111001111" => A <= "000000000000000000"; -- Line 125   Column 16   Coefficient 0.00000000
         when "011111010000" => A <= "000000000000000000"; -- Line 126   Column 1   Coefficient 0.00000000
         when "011111010001" => A <= "000000000000000000"; -- Line 126   Column 2   Coefficient 0.00000000
         when "011111010010" => A <= "000000001111000010"; -- Line 126   Column 3   Coefficient 0.00366974
         when "011111010011" => A <= "111110000010011110"; -- Line 126   Column 4   Coefficient -0.03064728
         when "011111010100" => A <= "010011010010100110"; -- Line 126   Column 5   Coefficient 0.30141449
         when "011111010101" => A <= "111101100111001110"; -- Line 126   Column 6   Coefficient -0.03730011
         when "011111010110" => A <= "000000110010101110"; -- Line 126   Column 7   Coefficient 0.01238251
         when "011111010111" => A <= "000000000001111110"; -- Line 126   Column 8   Coefficient 0.00048065
         when "011111011000" => A <= "000000000000000000"; -- Line 126   Column 9   Coefficient 0.00000000
         when "011111011001" => A <= "000000000000000000"; -- Line 126   Column 10   Coefficient 0.00000000
         when "011111011010" => A <= "000000000000000000"; -- Line 126   Column 11   Coefficient 0.00000000
         when "011111011011" => A <= "000000000000000000"; -- Line 126   Column 12   Coefficient 0.00000000
         when "011111011100" => A <= "000000000000000000"; -- Line 126   Column 13   Coefficient 0.00000000
         when "011111011101" => A <= "000000000000000000"; -- Line 126   Column 14   Coefficient 0.00000000
         when "011111011110" => A <= "000000000000000000"; -- Line 126   Column 15   Coefficient 0.00000000
         when "011111011111" => A <= "000000000000000000"; -- Line 126   Column 16   Coefficient 0.00000000
         when "011111100000" => A <= "000000000000000000"; -- Line 127   Column 1   Coefficient 0.00000000
         when "011111100001" => A <= "000000000000000000"; -- Line 127   Column 2   Coefficient 0.00000000
         when "011111100010" => A <= "000000010000011000"; -- Line 127   Column 3   Coefficient 0.00399780
         when "011111100011" => A <= "111101101011101110"; -- Line 127   Column 4   Coefficient -0.03620148
         when "011111100100" => A <= "010010110100110100"; -- Line 127   Column 5   Coefficient 0.29414368
         when "011111100101" => A <= "111110100000101100"; -- Line 127   Column 6   Coefficient -0.02326965
         when "011111100110" => A <= "000000101101010111"; -- Line 127   Column 7   Coefficient 0.01107407
         when "011111100111" => A <= "000000000001000010"; -- Line 127   Column 8   Coefficient 0.00025177
         when "011111101000" => A <= "000000000000000000"; -- Line 127   Column 9   Coefficient 0.00000000
         when "011111101001" => A <= "000000000000000000"; -- Line 127   Column 10   Coefficient 0.00000000
         when "011111101010" => A <= "000000000000000000"; -- Line 127   Column 11   Coefficient 0.00000000
         when "011111101011" => A <= "000000000000000000"; -- Line 127   Column 12   Coefficient 0.00000000
         when "011111101100" => A <= "000000000000000000"; -- Line 127   Column 13   Coefficient 0.00000000
         when "011111101101" => A <= "000000000000000000"; -- Line 127   Column 14   Coefficient 0.00000000
         when "011111101110" => A <= "000000000000000000"; -- Line 127   Column 15   Coefficient 0.00000000
         when "011111101111" => A <= "000000000000000000"; -- Line 127   Column 16   Coefficient 0.00000000
         when "011111110000" => A <= "000000000000000000"; -- Line 128   Column 1   Coefficient 0.00000000
         when "011111110001" => A <= "000000000000000000"; -- Line 128   Column 2   Coefficient 0.00000000
         when "011111110010" => A <= "000000001111111100"; -- Line 128   Column 3   Coefficient 0.00389099
         when "011111110011" => A <= "111101100000101101"; -- Line 128   Column 4   Coefficient -0.03889084
         when "011111110100" => A <= "010010000001100011"; -- Line 128   Column 5   Coefficient 0.28162766
         when "011111110101" => A <= "111111101010001000"; -- Line 128   Column 6   Coefficient -0.00534058
         when "011111110110" => A <= "000000100010100100"; -- Line 128   Column 7   Coefficient 0.00843811
         when "011111110111" => A <= "000000000001001000"; -- Line 128   Column 8   Coefficient 0.00027466
         when "011111111000" => A <= "000000000000000000"; -- Line 128   Column 9   Coefficient 0.00000000
         when "011111111001" => A <= "000000000000000000"; -- Line 128   Column 10   Coefficient 0.00000000
         when "011111111010" => A <= "000000000000000000"; -- Line 128   Column 11   Coefficient 0.00000000
         when "011111111011" => A <= "000000000000000000"; -- Line 128   Column 12   Coefficient 0.00000000
         when "011111111100" => A <= "000000000000000000"; -- Line 128   Column 13   Coefficient 0.00000000
         when "011111111101" => A <= "000000000000000000"; -- Line 128   Column 14   Coefficient 0.00000000
         when "011111111110" => A <= "000000000000000000"; -- Line 128   Column 15   Coefficient 0.00000000
         when "011111111111" => A <= "000000000000000000"; -- Line 128   Column 16   Coefficient 0.00000000
         when "100000000000" => A <= "000000000000000000"; -- Line 129   Column 1   Coefficient 0.00000000
         when "100000000001" => A <= "000000000000000000"; -- Line 129   Column 2   Coefficient 0.00000000
         when "100000000010" => A <= "000000001101001100"; -- Line 129   Column 3   Coefficient 0.00321960
         when "100000000011" => A <= "111101100010001110"; -- Line 129   Column 4   Coefficient -0.03852081
         when "100000000100" => A <= "010000111010100101"; -- Line 129   Column 5   Coefficient 0.26430130
         when "100000000101" => A <= "000000111110100110"; -- Line 129   Column 6   Coefficient 0.01528168
         when "100000000110" => A <= "000000010110010000"; -- Line 129   Column 7   Coefficient 0.00543213
         when "100000000111" => A <= "000000000001001011"; -- Line 129   Column 8   Coefficient 0.00028610
         when "100000001000" => A <= "000000000000000000"; -- Line 129   Column 9   Coefficient 0.00000000
         when "100000001001" => A <= "000000000000000000"; -- Line 129   Column 10   Coefficient 0.00000000
         when "100000001010" => A <= "000000000000000000"; -- Line 129   Column 11   Coefficient 0.00000000
         when "100000001011" => A <= "000000000000000000"; -- Line 129   Column 12   Coefficient 0.00000000
         when "100000001100" => A <= "000000000000000000"; -- Line 129   Column 13   Coefficient 0.00000000
         when "100000001101" => A <= "000000000000000000"; -- Line 129   Column 14   Coefficient 0.00000000
         when "100000001110" => A <= "000000000000000000"; -- Line 129   Column 15   Coefficient 0.00000000
         when "100000001111" => A <= "000000000000000000"; -- Line 129   Column 16   Coefficient 0.00000000
         when "100000010000" => A <= "000000000000000000"; -- Line 130   Column 1   Coefficient 0.00000000
         when "100000010001" => A <= "000000000000000000"; -- Line 130   Column 2   Coefficient 0.00000000
         when "100000010010" => A <= "000000001010110110"; -- Line 130   Column 3   Coefficient 0.00264740
         when "100000010011" => A <= "111101100010101111"; -- Line 130   Column 4   Coefficient -0.03839493
         when "100000010100" => A <= "001111111010100001"; -- Line 130   Column 5   Coefficient 0.24866104
         when "100000010101" => A <= "000010000100001011"; -- Line 130   Column 6   Coefficient 0.03226852
         when "100000010110" => A <= "000000010100110111"; -- Line 130   Column 7   Coefficient 0.00509262
         when "100000010111" => A <= "111111111110110111"; -- Line 130   Column 8   Coefficient -0.00027847
         when "100000011000" => A <= "000000000000000000"; -- Line 130   Column 9   Coefficient 0.00000000
         when "100000011001" => A <= "000000000000000000"; -- Line 130   Column 10   Coefficient 0.00000000
         when "100000011010" => A <= "000000000000000000"; -- Line 130   Column 11   Coefficient 0.00000000
         when "100000011011" => A <= "000000000000000000"; -- Line 130   Column 12   Coefficient 0.00000000
         when "100000011100" => A <= "000000000000000000"; -- Line 130   Column 13   Coefficient 0.00000000
         when "100000011101" => A <= "000000000000000000"; -- Line 130   Column 14   Coefficient 0.00000000
         when "100000011110" => A <= "000000000000000000"; -- Line 130   Column 15   Coefficient 0.00000000
         when "100000011111" => A <= "000000000000000000"; -- Line 130   Column 16   Coefficient 0.00000000
         when "100000100000" => A <= "000000000000000000"; -- Line 131   Column 1   Coefficient 0.00000000
         when "100000100001" => A <= "000000000000000000"; -- Line 131   Column 2   Coefficient 0.00000000
         when "100000100010" => A <= "000000001000010011"; -- Line 131   Column 3   Coefficient 0.00202560
         when "100000100011" => A <= "111101100110110000"; -- Line 131   Column 4   Coefficient -0.03741455
         when "100000100100" => A <= "001110110101010100"; -- Line 131   Column 5   Coefficient 0.23176575
         when "100000100101" => A <= "000011001010010011"; -- Line 131   Column 6   Coefficient 0.04938889
         when "100000100110" => A <= "000000010100111001"; -- Line 131   Column 7   Coefficient 0.00510025
         when "100000100111" => A <= "111111111100011110"; -- Line 131   Column 8   Coefficient -0.00086212
         when "100000101000" => A <= "111111111111111111"; -- Line 131   Column 9   Coefficient -0.00000381
         when "100000101001" => A <= "000000000000000000"; -- Line 131   Column 10   Coefficient 0.00000000
         when "100000101010" => A <= "000000000000000000"; -- Line 131   Column 11   Coefficient 0.00000000
         when "100000101011" => A <= "000000000000000000"; -- Line 131   Column 12   Coefficient 0.00000000
         when "100000101100" => A <= "000000000000000000"; -- Line 131   Column 13   Coefficient 0.00000000
         when "100000101101" => A <= "000000000000000000"; -- Line 131   Column 14   Coefficient 0.00000000
         when "100000101110" => A <= "000000000000000000"; -- Line 131   Column 15   Coefficient 0.00000000
         when "100000101111" => A <= "000000000000000000"; -- Line 131   Column 16   Coefficient 0.00000000
         when "100000110000" => A <= "000000000000000000"; -- Line 132   Column 1   Coefficient 0.00000000
         when "100000110001" => A <= "000000000000000000"; -- Line 132   Column 2   Coefficient 0.00000000
         when "100000110010" => A <= "000000000011111000"; -- Line 132   Column 3   Coefficient 0.00094604
         when "100000110011" => A <= "111101110100001010"; -- Line 132   Column 4   Coefficient -0.03414154
         when "100000110100" => A <= "001101100011111111"; -- Line 132   Column 5   Coefficient 0.21191025
         when "100000110101" => A <= "000100010011001101"; -- Line 132   Column 6   Coefficient 0.06718826
         when "100000110110" => A <= "000000010111101010"; -- Line 132   Column 7   Coefficient 0.00577545
         when "100000110111" => A <= "111111111001000110"; -- Line 132   Column 8   Coefficient -0.00168610
         when "100000111000" => A <= "000000000000000011"; -- Line 132   Column 9   Coefficient 0.00001144
         when "100000111001" => A <= "000000000000000000"; -- Line 132   Column 10   Coefficient 0.00000000
         when "100000111010" => A <= "000000000000000000"; -- Line 132   Column 11   Coefficient 0.00000000
         when "100000111011" => A <= "000000000000000000"; -- Line 132   Column 12   Coefficient 0.00000000
         when "100000111100" => A <= "000000000000000000"; -- Line 132   Column 13   Coefficient 0.00000000
         when "100000111101" => A <= "000000000000000000"; -- Line 132   Column 14   Coefficient 0.00000000
         when "100000111110" => A <= "000000000000000000"; -- Line 132   Column 15   Coefficient 0.00000000
         when "100000111111" => A <= "000000000000000000"; -- Line 132   Column 16   Coefficient 0.00000000
         when "100001000000" => A <= "000000000000000000"; -- Line 133   Column 1   Coefficient 0.00000000
         when "100001000001" => A <= "000000000000000000"; -- Line 133   Column 2   Coefficient 0.00000000
         when "100001000010" => A <= "111111111111010011"; -- Line 133   Column 3   Coefficient -0.00017166
         when "100001000011" => A <= "111110000101010011"; -- Line 133   Column 4   Coefficient -0.02995682
         when "100001000100" => A <= "001100001011101000"; -- Line 133   Column 5   Coefficient 0.19033813
         when "100001000101" => A <= "000101100000010101"; -- Line 133   Column 6   Coefficient 0.08601761
         when "100001000110" => A <= "000000011000110111"; -- Line 133   Column 7   Coefficient 0.00606918
         when "100001000111" => A <= "111111110110011111"; -- Line 133   Column 8   Coefficient -0.00232315
         when "100001001000" => A <= "000000000000000110"; -- Line 133   Column 9   Coefficient 0.00002289
         when "100001001001" => A <= "000000000000000000"; -- Line 133   Column 10   Coefficient 0.00000000
         when "100001001010" => A <= "000000000000000000"; -- Line 133   Column 11   Coefficient 0.00000000
         when "100001001011" => A <= "000000000000000000"; -- Line 133   Column 12   Coefficient 0.00000000
         when "100001001100" => A <= "000000000000000000"; -- Line 133   Column 13   Coefficient 0.00000000
         when "100001001101" => A <= "000000000000000000"; -- Line 133   Column 14   Coefficient 0.00000000
         when "100001001110" => A <= "000000000000000000"; -- Line 133   Column 15   Coefficient 0.00000000
         when "100001001111" => A <= "000000000000000000"; -- Line 133   Column 16   Coefficient 0.00000000
         when "100001010000" => A <= "000000000000000000"; -- Line 134   Column 1   Coefficient 0.00000000
         when "100001010001" => A <= "000000000000000000"; -- Line 134   Column 2   Coefficient 0.00000000
         when "100001010010" => A <= "111111111110010010"; -- Line 134   Column 3   Coefficient -0.00041962
         when "100001010011" => A <= "111110010000110000"; -- Line 134   Column 4   Coefficient -0.02716064
         when "100001010100" => A <= "001010101100000111"; -- Line 134   Column 5   Coefficient 0.16701889
         when "100001010101" => A <= "000111000101010101"; -- Line 134   Column 6   Coefficient 0.11067581
         when "100001010110" => A <= "000000000100100100"; -- Line 134   Column 7   Coefficient 0.00111389
         when "100001010111" => A <= "111111111010111001"; -- Line 134   Column 8   Coefficient -0.00124741
         when "100001011000" => A <= "000000000000000100"; -- Line 134   Column 9   Coefficient 0.00001526
         when "100001011001" => A <= "000000000000000000"; -- Line 134   Column 10   Coefficient 0.00000000
         when "100001011010" => A <= "000000000000000000"; -- Line 134   Column 11   Coefficient 0.00000000
         when "100001011011" => A <= "000000000000000000"; -- Line 134   Column 12   Coefficient 0.00000000
         when "100001011100" => A <= "000000000000000000"; -- Line 134   Column 13   Coefficient 0.00000000
         when "100001011101" => A <= "000000000000000000"; -- Line 134   Column 14   Coefficient 0.00000000
         when "100001011110" => A <= "000000000000000000"; -- Line 134   Column 15   Coefficient 0.00000000
         when "100001011111" => A <= "000000000000000000"; -- Line 134   Column 16   Coefficient 0.00000000
         when "100001100000" => A <= "000000000000000000"; -- Line 135   Column 1   Coefficient 0.00000000
         when "100001100001" => A <= "000000000000000000"; -- Line 135   Column 2   Coefficient 0.00000000
         when "100001100010" => A <= "111111111110100110"; -- Line 135   Column 3   Coefficient -0.00034332
         when "100001100011" => A <= "111110011011111010"; -- Line 135   Column 4   Coefficient -0.02443695
         when "100001100100" => A <= "001001000110101001"; -- Line 135   Column 5   Coefficient 0.14224625
         when "100001100101" => A <= "001000110101000000"; -- Line 135   Column 6   Coefficient 0.13793945
         when "100001100110" => A <= "111111100111100010"; -- Line 135   Column 7   Coefficient -0.00597382
         when "100001100111" => A <= "000000000010010011"; -- Line 135   Column 8   Coefficient 0.00056076
         when "100001101000" => A <= "000000000000000011"; -- Line 135   Column 9   Coefficient 0.00001144
         when "100001101001" => A <= "000000000000000000"; -- Line 135   Column 10   Coefficient 0.00000000
         when "100001101010" => A <= "000000000000000000"; -- Line 135   Column 11   Coefficient 0.00000000
         when "100001101011" => A <= "000000000000000000"; -- Line 135   Column 12   Coefficient 0.00000000
         when "100001101100" => A <= "000000000000000000"; -- Line 135   Column 13   Coefficient 0.00000000
         when "100001101101" => A <= "000000000000000000"; -- Line 135   Column 14   Coefficient 0.00000000
         when "100001101110" => A <= "000000000000000000"; -- Line 135   Column 15   Coefficient 0.00000000
         when "100001101111" => A <= "000000000000000000"; -- Line 135   Column 16   Coefficient 0.00000000
         when "100001110000" => A <= "000000000000000000"; -- Line 136   Column 1   Coefficient 0.00000000
         when "100001110001" => A <= "000000000000000000"; -- Line 136   Column 2   Coefficient 0.00000000
         when "100001110010" => A <= "111111111111001011"; -- Line 136   Column 3   Coefficient -0.00020218
         when "100001110011" => A <= "111110100110010011"; -- Line 136   Column 4   Coefficient -0.02190018
         when "100001110100" => A <= "000111100110110001"; -- Line 136   Column 5   Coefficient 0.11883926
         when "100001110101" => A <= "001010011001111000"; -- Line 136   Column 6   Coefficient 0.16256714
         when "100001110110" => A <= "111111010000101110"; -- Line 136   Column 7   Coefficient -0.01154327
         when "100001110111" => A <= "000000001001011000"; -- Line 136   Column 8   Coefficient 0.00228882
         when "100001111000" => A <= "111111111111110100"; -- Line 136   Column 9   Coefficient -0.00004578
         when "100001111001" => A <= "000000000000000000"; -- Line 136   Column 10   Coefficient 0.00000000
         when "100001111010" => A <= "000000000000000000"; -- Line 136   Column 11   Coefficient 0.00000000
         when "100001111011" => A <= "000000000000000000"; -- Line 136   Column 12   Coefficient 0.00000000
         when "100001111100" => A <= "000000000000000000"; -- Line 136   Column 13   Coefficient 0.00000000
         when "100001111101" => A <= "000000000000000000"; -- Line 136   Column 14   Coefficient 0.00000000
         when "100001111110" => A <= "000000000000000000"; -- Line 136   Column 15   Coefficient 0.00000000
         when "100001111111" => A <= "000000000000000000"; -- Line 136   Column 16   Coefficient 0.00000000
         when "100010000000" => A <= "000000000000000000"; -- Line 137   Column 1   Coefficient 0.00000000
         when "100010000001" => A <= "000000000000000000"; -- Line 137   Column 2   Coefficient 0.00000000
         when "100010000010" => A <= "000000000000000011"; -- Line 137   Column 3   Coefficient 0.00001144
         when "100010000011" => A <= "111110110001100001"; -- Line 137   Column 4   Coefficient -0.01916122
         when "100010000100" => A <= "000110000101110011"; -- Line 137   Column 5   Coefficient 0.09516525
         when "100010000101" => A <= "001011111101111010"; -- Line 137   Column 6   Coefficient 0.18698883
         when "100010000110" => A <= "111110111010000001"; -- Line 137   Column 7   Coefficient -0.01708603
         when "100010000111" => A <= "000000010001001000"; -- Line 137   Column 8   Coefficient 0.00418091
         when "100010001000" => A <= "111111111111100110"; -- Line 137   Column 9   Coefficient -0.00009918
         when "100010001001" => A <= "000000000000000000"; -- Line 137   Column 10   Coefficient 0.00000000
         when "100010001010" => A <= "000000000000000000"; -- Line 137   Column 11   Coefficient 0.00000000
         when "100010001011" => A <= "000000000000000000"; -- Line 137   Column 12   Coefficient 0.00000000
         when "100010001100" => A <= "000000000000000000"; -- Line 137   Column 13   Coefficient 0.00000000
         when "100010001101" => A <= "000000000000000000"; -- Line 137   Column 14   Coefficient 0.00000000
         when "100010001110" => A <= "000000000000000000"; -- Line 137   Column 15   Coefficient 0.00000000
         when "100010001111" => A <= "000000000000000000"; -- Line 137   Column 16   Coefficient 0.00000000
         when "100010010000" => A <= "000000000000000000"; -- Line 138   Column 1   Coefficient 0.00000000
         when "100010010001" => A <= "000000000000000000"; -- Line 138   Column 2   Coefficient 0.00000000
         when "100010010010" => A <= "000000000000001001"; -- Line 138   Column 3   Coefficient 0.00003433
         when "100010010011" => A <= "111111000100111001"; -- Line 138   Column 4   Coefficient -0.01443100
         when "100010010100" => A <= "000100010010000101"; -- Line 138   Column 5   Coefficient 0.06691360
         when "100010010101" => A <= "001101110100101001"; -- Line 138   Column 6   Coefficient 0.21597672
         when "100010010110" => A <= "111110011010010101"; -- Line 138   Column 7   Coefficient -0.02482224
         when "100010010111" => A <= "000000011001110100"; -- Line 138   Column 8   Coefficient 0.00630188
         when "100010011000" => A <= "000000000000000111"; -- Line 138   Column 9   Coefficient 0.00002670
         when "100010011001" => A <= "000000000000000000"; -- Line 138   Column 10   Coefficient 0.00000000
         when "100010011010" => A <= "000000000000000000"; -- Line 138   Column 11   Coefficient 0.00000000
         when "100010011011" => A <= "000000000000000000"; -- Line 138   Column 12   Coefficient 0.00000000
         when "100010011100" => A <= "000000000000000000"; -- Line 138   Column 13   Coefficient 0.00000000
         when "100010011101" => A <= "000000000000000000"; -- Line 138   Column 14   Coefficient 0.00000000
         when "100010011110" => A <= "000000000000000000"; -- Line 138   Column 15   Coefficient 0.00000000
         when "100010011111" => A <= "000000000000000000"; -- Line 138   Column 16   Coefficient 0.00000000
         when "100010100000" => A <= "000000000000000000"; -- Line 139   Column 1   Coefficient 0.00000000
         when "100010100001" => A <= "000000000000000000"; -- Line 139   Column 2   Coefficient 0.00000000
         when "100010100010" => A <= "000000000000000000"; -- Line 139   Column 3   Coefficient 0.00000000
         when "100010100011" => A <= "111111011001111001"; -- Line 139   Column 4   Coefficient -0.00930405
         when "100010100100" => A <= "000010011110111100"; -- Line 139   Column 5   Coefficient 0.03880310
         when "100010100101" => A <= "001111100101110011"; -- Line 139   Column 6   Coefficient 0.24360275
         when "100010100110" => A <= "111101111110110001"; -- Line 139   Column 7   Coefficient -0.03155136
         when "100010100111" => A <= "000000100001110011"; -- Line 139   Column 8   Coefficient 0.00825119
         when "100010101000" => A <= "000000000000110011"; -- Line 139   Column 9   Coefficient 0.00019455
         when "100010101001" => A <= "000000000000000000"; -- Line 139   Column 10   Coefficient 0.00000000
         when "100010101010" => A <= "000000000000000000"; -- Line 139   Column 11   Coefficient 0.00000000
         when "100010101011" => A <= "000000000000000000"; -- Line 139   Column 12   Coefficient 0.00000000
         when "100010101100" => A <= "000000000000000000"; -- Line 139   Column 13   Coefficient 0.00000000
         when "100010101101" => A <= "000000000000000000"; -- Line 139   Column 14   Coefficient 0.00000000
         when "100010101110" => A <= "000000000000000000"; -- Line 139   Column 15   Coefficient 0.00000000
         when "100010101111" => A <= "000000000000000000"; -- Line 139   Column 16   Coefficient 0.00000000
         when "100010110000" => A <= "000000000000000000"; -- Line 140   Column 1   Coefficient 0.00000000
         when "100010110001" => A <= "000000000000000000"; -- Line 140   Column 2   Coefficient 0.00000000
         when "100010110010" => A <= "000000000000000000"; -- Line 140   Column 3   Coefficient 0.00000000
         when "100010110011" => A <= "111111110001010101"; -- Line 140   Column 4   Coefficient -0.00358200
         when "100010110100" => A <= "000000100101011001"; -- Line 140   Column 5   Coefficient 0.00912857
         when "100010110101" => A <= "010001011110001011"; -- Line 140   Column 6   Coefficient 0.27299118
         when "100010110110" => A <= "111101011101101101"; -- Line 140   Column 7   Coefficient -0.03962326
         when "100010110111" => A <= "000000101011110101"; -- Line 140   Column 8   Coefficient 0.01070023
         when "100010111000" => A <= "000000000001100101"; -- Line 140   Column 9   Coefficient 0.00038528
         when "100010111001" => A <= "000000000000000000"; -- Line 140   Column 10   Coefficient 0.00000000
         when "100010111010" => A <= "000000000000000000"; -- Line 140   Column 11   Coefficient 0.00000000
         when "100010111011" => A <= "000000000000000000"; -- Line 140   Column 12   Coefficient 0.00000000
         when "100010111100" => A <= "000000000000000000"; -- Line 140   Column 13   Coefficient 0.00000000
         when "100010111101" => A <= "000000000000000000"; -- Line 140   Column 14   Coefficient 0.00000000
         when "100010111110" => A <= "000000000000000000"; -- Line 140   Column 15   Coefficient 0.00000000
         when "100010111111" => A <= "000000000000000000"; -- Line 140   Column 16   Coefficient 0.00000000
         when "100011000000" => A <= "000000000000000000"; -- Line 141   Column 1   Coefficient 0.00000000
         when "100011000001" => A <= "000000000000000000"; -- Line 141   Column 2   Coefficient 0.00000000
         when "100011000010" => A <= "000000000000000000"; -- Line 141   Column 3   Coefficient 0.00000000
         when "100011000011" => A <= "000000000111011010"; -- Line 141   Column 4   Coefficient 0.00180817
         when "100011000100" => A <= "111110110101100100"; -- Line 141   Column 5   Coefficient -0.01817322
         when "100011000101" => A <= "010011000101100111"; -- Line 141   Column 6   Coefficient 0.29824448
         when "100011000110" => A <= "111101000110110001"; -- Line 141   Column 7   Coefficient -0.04522324
         when "100011000111" => A <= "000000110100010110"; -- Line 141   Column 8   Coefficient 0.01277924
         when "100011001000" => A <= "000000000010010101"; -- Line 141   Column 9   Coefficient 0.00056839
         when "100011001001" => A <= "000000000000000000"; -- Line 141   Column 10   Coefficient 0.00000000
         when "100011001010" => A <= "000000000000000000"; -- Line 141   Column 11   Coefficient 0.00000000
         when "100011001011" => A <= "000000000000000000"; -- Line 141   Column 12   Coefficient 0.00000000
         when "100011001100" => A <= "000000000000000000"; -- Line 141   Column 13   Coefficient 0.00000000
         when "100011001101" => A <= "000000000000000000"; -- Line 141   Column 14   Coefficient 0.00000000
         when "100011001110" => A <= "000000000000000000"; -- Line 141   Column 15   Coefficient 0.00000000
         when "100011001111" => A <= "000000000000000000"; -- Line 141   Column 16   Coefficient 0.00000000
         when "100011010000" => A <= "000000000000000000"; -- Line 142   Column 1   Coefficient 0.00000000
         when "100011010001" => A <= "000000000000000000"; -- Line 142   Column 2   Coefficient 0.00000000
         when "100011010010" => A <= "000000000000000000"; -- Line 142   Column 3   Coefficient 0.00000000
         when "100011010011" => A <= "000000001111000010"; -- Line 142   Column 4   Coefficient 0.00366974
         when "100011010100" => A <= "111110000010011110"; -- Line 142   Column 5   Coefficient -0.03064728
         when "100011010101" => A <= "010011010010100110"; -- Line 142   Column 6   Coefficient 0.30141449
         when "100011010110" => A <= "111101100111001110"; -- Line 142   Column 7   Coefficient -0.03730011
         when "100011010111" => A <= "000000110010101110"; -- Line 142   Column 8   Coefficient 0.01238251
         when "100011011000" => A <= "000000000001111110"; -- Line 142   Column 9   Coefficient 0.00048065
         when "100011011001" => A <= "000000000000000000"; -- Line 142   Column 10   Coefficient 0.00000000
         when "100011011010" => A <= "000000000000000000"; -- Line 142   Column 11   Coefficient 0.00000000
         when "100011011011" => A <= "000000000000000000"; -- Line 142   Column 12   Coefficient 0.00000000
         when "100011011100" => A <= "000000000000000000"; -- Line 142   Column 13   Coefficient 0.00000000
         when "100011011101" => A <= "000000000000000000"; -- Line 142   Column 14   Coefficient 0.00000000
         when "100011011110" => A <= "000000000000000000"; -- Line 142   Column 15   Coefficient 0.00000000
         when "100011011111" => A <= "000000000000000000"; -- Line 142   Column 16   Coefficient 0.00000000
         when "100011100000" => A <= "000000000000000000"; -- Line 143   Column 1   Coefficient 0.00000000
         when "100011100001" => A <= "000000000000000000"; -- Line 143   Column 2   Coefficient 0.00000000
         when "100011100010" => A <= "000000000000000000"; -- Line 143   Column 3   Coefficient 0.00000000
         when "100011100011" => A <= "000000010000011000"; -- Line 143   Column 4   Coefficient 0.00399780
         when "100011100100" => A <= "111101101011101110"; -- Line 143   Column 5   Coefficient -0.03620148
         when "100011100101" => A <= "010010110100110100"; -- Line 143   Column 6   Coefficient 0.29414368
         when "100011100110" => A <= "111110100000101100"; -- Line 143   Column 7   Coefficient -0.02326965
         when "100011100111" => A <= "000000101101010111"; -- Line 143   Column 8   Coefficient 0.01107407
         when "100011101000" => A <= "000000000001000010"; -- Line 143   Column 9   Coefficient 0.00025177
         when "100011101001" => A <= "000000000000000000"; -- Line 143   Column 10   Coefficient 0.00000000
         when "100011101010" => A <= "000000000000000000"; -- Line 143   Column 11   Coefficient 0.00000000
         when "100011101011" => A <= "000000000000000000"; -- Line 143   Column 12   Coefficient 0.00000000
         when "100011101100" => A <= "000000000000000000"; -- Line 143   Column 13   Coefficient 0.00000000
         when "100011101101" => A <= "000000000000000000"; -- Line 143   Column 14   Coefficient 0.00000000
         when "100011101110" => A <= "000000000000000000"; -- Line 143   Column 15   Coefficient 0.00000000
         when "100011101111" => A <= "000000000000000000"; -- Line 143   Column 16   Coefficient 0.00000000
         when "100011110000" => A <= "000000000000000000"; -- Line 144   Column 1   Coefficient 0.00000000
         when "100011110001" => A <= "000000000000000000"; -- Line 144   Column 2   Coefficient 0.00000000
         when "100011110010" => A <= "000000000000000000"; -- Line 144   Column 3   Coefficient 0.00000000
         when "100011110011" => A <= "000000001111111100"; -- Line 144   Column 4   Coefficient 0.00389099
         when "100011110100" => A <= "111101100000101101"; -- Line 144   Column 5   Coefficient -0.03889084
         when "100011110101" => A <= "010010000001100011"; -- Line 144   Column 6   Coefficient 0.28162766
         when "100011110110" => A <= "111111101010001000"; -- Line 144   Column 7   Coefficient -0.00534058
         when "100011110111" => A <= "000000100010100100"; -- Line 144   Column 8   Coefficient 0.00843811
         when "100011111000" => A <= "000000000001001000"; -- Line 144   Column 9   Coefficient 0.00027466
         when "100011111001" => A <= "000000000000000000"; -- Line 144   Column 10   Coefficient 0.00000000
         when "100011111010" => A <= "000000000000000000"; -- Line 144   Column 11   Coefficient 0.00000000
         when "100011111011" => A <= "000000000000000000"; -- Line 144   Column 12   Coefficient 0.00000000
         when "100011111100" => A <= "000000000000000000"; -- Line 144   Column 13   Coefficient 0.00000000
         when "100011111101" => A <= "000000000000000000"; -- Line 144   Column 14   Coefficient 0.00000000
         when "100011111110" => A <= "000000000000000000"; -- Line 144   Column 15   Coefficient 0.00000000
         when "100011111111" => A <= "000000000000000000"; -- Line 144   Column 16   Coefficient 0.00000000
         when "100100000000" => A <= "000000000000000000"; -- Line 145   Column 1   Coefficient 0.00000000
         when "100100000001" => A <= "000000000000000000"; -- Line 145   Column 2   Coefficient 0.00000000
         when "100100000010" => A <= "000000000000000000"; -- Line 145   Column 3   Coefficient 0.00000000
         when "100100000011" => A <= "000000001101001100"; -- Line 145   Column 4   Coefficient 0.00321960
         when "100100000100" => A <= "111101100010001110"; -- Line 145   Column 5   Coefficient -0.03852081
         when "100100000101" => A <= "010000111010100101"; -- Line 145   Column 6   Coefficient 0.26430130
         when "100100000110" => A <= "000000111110100110"; -- Line 145   Column 7   Coefficient 0.01528168
         when "100100000111" => A <= "000000010110010000"; -- Line 145   Column 8   Coefficient 0.00543213
         when "100100001000" => A <= "000000000001001011"; -- Line 145   Column 9   Coefficient 0.00028610
         when "100100001001" => A <= "000000000000000000"; -- Line 145   Column 10   Coefficient 0.00000000
         when "100100001010" => A <= "000000000000000000"; -- Line 145   Column 11   Coefficient 0.00000000
         when "100100001011" => A <= "000000000000000000"; -- Line 145   Column 12   Coefficient 0.00000000
         when "100100001100" => A <= "000000000000000000"; -- Line 145   Column 13   Coefficient 0.00000000
         when "100100001101" => A <= "000000000000000000"; -- Line 145   Column 14   Coefficient 0.00000000
         when "100100001110" => A <= "000000000000000000"; -- Line 145   Column 15   Coefficient 0.00000000
         when "100100001111" => A <= "000000000000000000"; -- Line 145   Column 16   Coefficient 0.00000000
         when "100100010000" => A <= "000000000000000000"; -- Line 146   Column 1   Coefficient 0.00000000
         when "100100010001" => A <= "000000000000000000"; -- Line 146   Column 2   Coefficient 0.00000000
         when "100100010010" => A <= "000000000000000000"; -- Line 146   Column 3   Coefficient 0.00000000
         when "100100010011" => A <= "000000001010110110"; -- Line 146   Column 4   Coefficient 0.00264740
         when "100100010100" => A <= "111101100010101111"; -- Line 146   Column 5   Coefficient -0.03839493
         when "100100010101" => A <= "001111111010100001"; -- Line 146   Column 6   Coefficient 0.24866104
         when "100100010110" => A <= "000010000100001011"; -- Line 146   Column 7   Coefficient 0.03226852
         when "100100010111" => A <= "000000010100110111"; -- Line 146   Column 8   Coefficient 0.00509262
         when "100100011000" => A <= "111111111110110111"; -- Line 146   Column 9   Coefficient -0.00027847
         when "100100011001" => A <= "000000000000000000"; -- Line 146   Column 10   Coefficient 0.00000000
         when "100100011010" => A <= "000000000000000000"; -- Line 146   Column 11   Coefficient 0.00000000
         when "100100011011" => A <= "000000000000000000"; -- Line 146   Column 12   Coefficient 0.00000000
         when "100100011100" => A <= "000000000000000000"; -- Line 146   Column 13   Coefficient 0.00000000
         when "100100011101" => A <= "000000000000000000"; -- Line 146   Column 14   Coefficient 0.00000000
         when "100100011110" => A <= "000000000000000000"; -- Line 146   Column 15   Coefficient 0.00000000
         when "100100011111" => A <= "000000000000000000"; -- Line 146   Column 16   Coefficient 0.00000000
         when "100100100000" => A <= "000000000000000000"; -- Line 147   Column 1   Coefficient 0.00000000
         when "100100100001" => A <= "000000000000000000"; -- Line 147   Column 2   Coefficient 0.00000000
         when "100100100010" => A <= "000000000000000000"; -- Line 147   Column 3   Coefficient 0.00000000
         when "100100100011" => A <= "000000001000010011"; -- Line 147   Column 4   Coefficient 0.00202560
         when "100100100100" => A <= "111101100110110000"; -- Line 147   Column 5   Coefficient -0.03741455
         when "100100100101" => A <= "001110110101010100"; -- Line 147   Column 6   Coefficient 0.23176575
         when "100100100110" => A <= "000011001010010011"; -- Line 147   Column 7   Coefficient 0.04938889
         when "100100100111" => A <= "000000010100111001"; -- Line 147   Column 8   Coefficient 0.00510025
         when "100100101000" => A <= "111111111100011110"; -- Line 147   Column 9   Coefficient -0.00086212
         when "100100101001" => A <= "111111111111111111"; -- Line 147   Column 10   Coefficient -0.00000381
         when "100100101010" => A <= "000000000000000000"; -- Line 147   Column 11   Coefficient 0.00000000
         when "100100101011" => A <= "000000000000000000"; -- Line 147   Column 12   Coefficient 0.00000000
         when "100100101100" => A <= "000000000000000000"; -- Line 147   Column 13   Coefficient 0.00000000
         when "100100101101" => A <= "000000000000000000"; -- Line 147   Column 14   Coefficient 0.00000000
         when "100100101110" => A <= "000000000000000000"; -- Line 147   Column 15   Coefficient 0.00000000
         when "100100101111" => A <= "000000000000000000"; -- Line 147   Column 16   Coefficient 0.00000000
         when "100100110000" => A <= "000000000000000000"; -- Line 148   Column 1   Coefficient 0.00000000
         when "100100110001" => A <= "000000000000000000"; -- Line 148   Column 2   Coefficient 0.00000000
         when "100100110010" => A <= "000000000000000000"; -- Line 148   Column 3   Coefficient 0.00000000
         when "100100110011" => A <= "000000000011111000"; -- Line 148   Column 4   Coefficient 0.00094604
         when "100100110100" => A <= "111101110100001010"; -- Line 148   Column 5   Coefficient -0.03414154
         when "100100110101" => A <= "001101100011111111"; -- Line 148   Column 6   Coefficient 0.21191025
         when "100100110110" => A <= "000100010011001101"; -- Line 148   Column 7   Coefficient 0.06718826
         when "100100110111" => A <= "000000010111101010"; -- Line 148   Column 8   Coefficient 0.00577545
         when "100100111000" => A <= "111111111001000110"; -- Line 148   Column 9   Coefficient -0.00168610
         when "100100111001" => A <= "000000000000000011"; -- Line 148   Column 10   Coefficient 0.00001144
         when "100100111010" => A <= "000000000000000000"; -- Line 148   Column 11   Coefficient 0.00000000
         when "100100111011" => A <= "000000000000000000"; -- Line 148   Column 12   Coefficient 0.00000000
         when "100100111100" => A <= "000000000000000000"; -- Line 148   Column 13   Coefficient 0.00000000
         when "100100111101" => A <= "000000000000000000"; -- Line 148   Column 14   Coefficient 0.00000000
         when "100100111110" => A <= "000000000000000000"; -- Line 148   Column 15   Coefficient 0.00000000
         when "100100111111" => A <= "000000000000000000"; -- Line 148   Column 16   Coefficient 0.00000000
         when "100101000000" => A <= "000000000000000000"; -- Line 149   Column 1   Coefficient 0.00000000
         when "100101000001" => A <= "000000000000000000"; -- Line 149   Column 2   Coefficient 0.00000000
         when "100101000010" => A <= "000000000000000000"; -- Line 149   Column 3   Coefficient 0.00000000
         when "100101000011" => A <= "111111111111010011"; -- Line 149   Column 4   Coefficient -0.00017166
         when "100101000100" => A <= "111110000101010011"; -- Line 149   Column 5   Coefficient -0.02995682
         when "100101000101" => A <= "001100001011101000"; -- Line 149   Column 6   Coefficient 0.19033813
         when "100101000110" => A <= "000101100000010101"; -- Line 149   Column 7   Coefficient 0.08601761
         when "100101000111" => A <= "000000011000110111"; -- Line 149   Column 8   Coefficient 0.00606918
         when "100101001000" => A <= "111111110110011111"; -- Line 149   Column 9   Coefficient -0.00232315
         when "100101001001" => A <= "000000000000000110"; -- Line 149   Column 10   Coefficient 0.00002289
         when "100101001010" => A <= "000000000000000000"; -- Line 149   Column 11   Coefficient 0.00000000
         when "100101001011" => A <= "000000000000000000"; -- Line 149   Column 12   Coefficient 0.00000000
         when "100101001100" => A <= "000000000000000000"; -- Line 149   Column 13   Coefficient 0.00000000
         when "100101001101" => A <= "000000000000000000"; -- Line 149   Column 14   Coefficient 0.00000000
         when "100101001110" => A <= "000000000000000000"; -- Line 149   Column 15   Coefficient 0.00000000
         when "100101001111" => A <= "000000000000000000"; -- Line 149   Column 16   Coefficient 0.00000000
         when "100101010000" => A <= "000000000000000000"; -- Line 150   Column 1   Coefficient 0.00000000
         when "100101010001" => A <= "000000000000000000"; -- Line 150   Column 2   Coefficient 0.00000000
         when "100101010010" => A <= "000000000000000000"; -- Line 150   Column 3   Coefficient 0.00000000
         when "100101010011" => A <= "111111111110010010"; -- Line 150   Column 4   Coefficient -0.00041962
         when "100101010100" => A <= "111110010000110000"; -- Line 150   Column 5   Coefficient -0.02716064
         when "100101010101" => A <= "001010101100000111"; -- Line 150   Column 6   Coefficient 0.16701889
         when "100101010110" => A <= "000111000101010101"; -- Line 150   Column 7   Coefficient 0.11067581
         when "100101010111" => A <= "000000000100100100"; -- Line 150   Column 8   Coefficient 0.00111389
         when "100101011000" => A <= "111111111010111001"; -- Line 150   Column 9   Coefficient -0.00124741
         when "100101011001" => A <= "000000000000000100"; -- Line 150   Column 10   Coefficient 0.00001526
         when "100101011010" => A <= "000000000000000000"; -- Line 150   Column 11   Coefficient 0.00000000
         when "100101011011" => A <= "000000000000000000"; -- Line 150   Column 12   Coefficient 0.00000000
         when "100101011100" => A <= "000000000000000000"; -- Line 150   Column 13   Coefficient 0.00000000
         when "100101011101" => A <= "000000000000000000"; -- Line 150   Column 14   Coefficient 0.00000000
         when "100101011110" => A <= "000000000000000000"; -- Line 150   Column 15   Coefficient 0.00000000
         when "100101011111" => A <= "000000000000000000"; -- Line 150   Column 16   Coefficient 0.00000000
         when "100101100000" => A <= "000000000000000000"; -- Line 151   Column 1   Coefficient 0.00000000
         when "100101100001" => A <= "000000000000000000"; -- Line 151   Column 2   Coefficient 0.00000000
         when "100101100010" => A <= "000000000000000000"; -- Line 151   Column 3   Coefficient 0.00000000
         when "100101100011" => A <= "111111111110100110"; -- Line 151   Column 4   Coefficient -0.00034332
         when "100101100100" => A <= "111110011011111010"; -- Line 151   Column 5   Coefficient -0.02443695
         when "100101100101" => A <= "001001000110101001"; -- Line 151   Column 6   Coefficient 0.14224625
         when "100101100110" => A <= "001000110101000000"; -- Line 151   Column 7   Coefficient 0.13793945
         when "100101100111" => A <= "111111100111100010"; -- Line 151   Column 8   Coefficient -0.00597382
         when "100101101000" => A <= "000000000010010011"; -- Line 151   Column 9   Coefficient 0.00056076
         when "100101101001" => A <= "000000000000000011"; -- Line 151   Column 10   Coefficient 0.00001144
         when "100101101010" => A <= "000000000000000000"; -- Line 151   Column 11   Coefficient 0.00000000
         when "100101101011" => A <= "000000000000000000"; -- Line 151   Column 12   Coefficient 0.00000000
         when "100101101100" => A <= "000000000000000000"; -- Line 151   Column 13   Coefficient 0.00000000
         when "100101101101" => A <= "000000000000000000"; -- Line 151   Column 14   Coefficient 0.00000000
         when "100101101110" => A <= "000000000000000000"; -- Line 151   Column 15   Coefficient 0.00000000
         when "100101101111" => A <= "000000000000000000"; -- Line 151   Column 16   Coefficient 0.00000000
         when "100101110000" => A <= "000000000000000000"; -- Line 152   Column 1   Coefficient 0.00000000
         when "100101110001" => A <= "000000000000000000"; -- Line 152   Column 2   Coefficient 0.00000000
         when "100101110010" => A <= "000000000000000000"; -- Line 152   Column 3   Coefficient 0.00000000
         when "100101110011" => A <= "111111111111001011"; -- Line 152   Column 4   Coefficient -0.00020218
         when "100101110100" => A <= "111110100110010011"; -- Line 152   Column 5   Coefficient -0.02190018
         when "100101110101" => A <= "000111100110110001"; -- Line 152   Column 6   Coefficient 0.11883926
         when "100101110110" => A <= "001010011001111000"; -- Line 152   Column 7   Coefficient 0.16256714
         when "100101110111" => A <= "111111010000101110"; -- Line 152   Column 8   Coefficient -0.01154327
         when "100101111000" => A <= "000000001001011000"; -- Line 152   Column 9   Coefficient 0.00228882
         when "100101111001" => A <= "111111111111110100"; -- Line 152   Column 10   Coefficient -0.00004578
         when "100101111010" => A <= "000000000000000000"; -- Line 152   Column 11   Coefficient 0.00000000
         when "100101111011" => A <= "000000000000000000"; -- Line 152   Column 12   Coefficient 0.00000000
         when "100101111100" => A <= "000000000000000000"; -- Line 152   Column 13   Coefficient 0.00000000
         when "100101111101" => A <= "000000000000000000"; -- Line 152   Column 14   Coefficient 0.00000000
         when "100101111110" => A <= "000000000000000000"; -- Line 152   Column 15   Coefficient 0.00000000
         when "100101111111" => A <= "000000000000000000"; -- Line 152   Column 16   Coefficient 0.00000000
         when "100110000000" => A <= "000000000000000000"; -- Line 153   Column 1   Coefficient 0.00000000
         when "100110000001" => A <= "000000000000000000"; -- Line 153   Column 2   Coefficient 0.00000000
         when "100110000010" => A <= "000000000000000000"; -- Line 153   Column 3   Coefficient 0.00000000
         when "100110000011" => A <= "000000000000000011"; -- Line 153   Column 4   Coefficient 0.00001144
         when "100110000100" => A <= "111110110001100001"; -- Line 153   Column 5   Coefficient -0.01916122
         when "100110000101" => A <= "000110000101110011"; -- Line 153   Column 6   Coefficient 0.09516525
         when "100110000110" => A <= "001011111101111010"; -- Line 153   Column 7   Coefficient 0.18698883
         when "100110000111" => A <= "111110111010000001"; -- Line 153   Column 8   Coefficient -0.01708603
         when "100110001000" => A <= "000000010001001000"; -- Line 153   Column 9   Coefficient 0.00418091
         when "100110001001" => A <= "111111111111100110"; -- Line 153   Column 10   Coefficient -0.00009918
         when "100110001010" => A <= "000000000000000000"; -- Line 153   Column 11   Coefficient 0.00000000
         when "100110001011" => A <= "000000000000000000"; -- Line 153   Column 12   Coefficient 0.00000000
         when "100110001100" => A <= "000000000000000000"; -- Line 153   Column 13   Coefficient 0.00000000
         when "100110001101" => A <= "000000000000000000"; -- Line 153   Column 14   Coefficient 0.00000000
         when "100110001110" => A <= "000000000000000000"; -- Line 153   Column 15   Coefficient 0.00000000
         when "100110001111" => A <= "000000000000000000"; -- Line 153   Column 16   Coefficient 0.00000000
         when "100110010000" => A <= "000000000000000000"; -- Line 154   Column 1   Coefficient 0.00000000
         when "100110010001" => A <= "000000000000000000"; -- Line 154   Column 2   Coefficient 0.00000000
         when "100110010010" => A <= "000000000000000000"; -- Line 154   Column 3   Coefficient 0.00000000
         when "100110010011" => A <= "000000000000001001"; -- Line 154   Column 4   Coefficient 0.00003433
         when "100110010100" => A <= "111111000100111001"; -- Line 154   Column 5   Coefficient -0.01443100
         when "100110010101" => A <= "000100010010000101"; -- Line 154   Column 6   Coefficient 0.06691360
         when "100110010110" => A <= "001101110100101001"; -- Line 154   Column 7   Coefficient 0.21597672
         when "100110010111" => A <= "111110011010010101"; -- Line 154   Column 8   Coefficient -0.02482224
         when "100110011000" => A <= "000000011001110100"; -- Line 154   Column 9   Coefficient 0.00630188
         when "100110011001" => A <= "000000000000000111"; -- Line 154   Column 10   Coefficient 0.00002670
         when "100110011010" => A <= "000000000000000000"; -- Line 154   Column 11   Coefficient 0.00000000
         when "100110011011" => A <= "000000000000000000"; -- Line 154   Column 12   Coefficient 0.00000000
         when "100110011100" => A <= "000000000000000000"; -- Line 154   Column 13   Coefficient 0.00000000
         when "100110011101" => A <= "000000000000000000"; -- Line 154   Column 14   Coefficient 0.00000000
         when "100110011110" => A <= "000000000000000000"; -- Line 154   Column 15   Coefficient 0.00000000
         when "100110011111" => A <= "000000000000000000"; -- Line 154   Column 16   Coefficient 0.00000000
         when "100110100000" => A <= "000000000000000000"; -- Line 155   Column 1   Coefficient 0.00000000
         when "100110100001" => A <= "000000000000000000"; -- Line 155   Column 2   Coefficient 0.00000000
         when "100110100010" => A <= "000000000000000000"; -- Line 155   Column 3   Coefficient 0.00000000
         when "100110100011" => A <= "000000000000000000"; -- Line 155   Column 4   Coefficient 0.00000000
         when "100110100100" => A <= "111111011001111001"; -- Line 155   Column 5   Coefficient -0.00930405
         when "100110100101" => A <= "000010011110111100"; -- Line 155   Column 6   Coefficient 0.03880310
         when "100110100110" => A <= "001111100101110011"; -- Line 155   Column 7   Coefficient 0.24360275
         when "100110100111" => A <= "111101111110110001"; -- Line 155   Column 8   Coefficient -0.03155136
         when "100110101000" => A <= "000000100001110011"; -- Line 155   Column 9   Coefficient 0.00825119
         when "100110101001" => A <= "000000000000110011"; -- Line 155   Column 10   Coefficient 0.00019455
         when "100110101010" => A <= "000000000000000000"; -- Line 155   Column 11   Coefficient 0.00000000
         when "100110101011" => A <= "000000000000000000"; -- Line 155   Column 12   Coefficient 0.00000000
         when "100110101100" => A <= "000000000000000000"; -- Line 155   Column 13   Coefficient 0.00000000
         when "100110101101" => A <= "000000000000000000"; -- Line 155   Column 14   Coefficient 0.00000000
         when "100110101110" => A <= "000000000000000000"; -- Line 155   Column 15   Coefficient 0.00000000
         when "100110101111" => A <= "000000000000000000"; -- Line 155   Column 16   Coefficient 0.00000000
         when "100110110000" => A <= "000000000000000000"; -- Line 156   Column 1   Coefficient 0.00000000
         when "100110110001" => A <= "000000000000000000"; -- Line 156   Column 2   Coefficient 0.00000000
         when "100110110010" => A <= "000000000000000000"; -- Line 156   Column 3   Coefficient 0.00000000
         when "100110110011" => A <= "000000000000000000"; -- Line 156   Column 4   Coefficient 0.00000000
         when "100110110100" => A <= "111111110001010101"; -- Line 156   Column 5   Coefficient -0.00358200
         when "100110110101" => A <= "000000100101011001"; -- Line 156   Column 6   Coefficient 0.00912857
         when "100110110110" => A <= "010001011110001011"; -- Line 156   Column 7   Coefficient 0.27299118
         when "100110110111" => A <= "111101011101101101"; -- Line 156   Column 8   Coefficient -0.03962326
         when "100110111000" => A <= "000000101011110101"; -- Line 156   Column 9   Coefficient 0.01070023
         when "100110111001" => A <= "000000000001100101"; -- Line 156   Column 10   Coefficient 0.00038528
         when "100110111010" => A <= "000000000000000000"; -- Line 156   Column 11   Coefficient 0.00000000
         when "100110111011" => A <= "000000000000000000"; -- Line 156   Column 12   Coefficient 0.00000000
         when "100110111100" => A <= "000000000000000000"; -- Line 156   Column 13   Coefficient 0.00000000
         when "100110111101" => A <= "000000000000000000"; -- Line 156   Column 14   Coefficient 0.00000000
         when "100110111110" => A <= "000000000000000000"; -- Line 156   Column 15   Coefficient 0.00000000
         when "100110111111" => A <= "000000000000000000"; -- Line 156   Column 16   Coefficient 0.00000000
         when "100111000000" => A <= "000000000000000000"; -- Line 157   Column 1   Coefficient 0.00000000
         when "100111000001" => A <= "000000000000000000"; -- Line 157   Column 2   Coefficient 0.00000000
         when "100111000010" => A <= "000000000000000000"; -- Line 157   Column 3   Coefficient 0.00000000
         when "100111000011" => A <= "000000000000000000"; -- Line 157   Column 4   Coefficient 0.00000000
         when "100111000100" => A <= "000000000111011010"; -- Line 157   Column 5   Coefficient 0.00180817
         when "100111000101" => A <= "111110110101100100"; -- Line 157   Column 6   Coefficient -0.01817322
         when "100111000110" => A <= "010011000101100111"; -- Line 157   Column 7   Coefficient 0.29824448
         when "100111000111" => A <= "111101000110110001"; -- Line 157   Column 8   Coefficient -0.04522324
         when "100111001000" => A <= "000000110100010110"; -- Line 157   Column 9   Coefficient 0.01277924
         when "100111001001" => A <= "000000000010010101"; -- Line 157   Column 10   Coefficient 0.00056839
         when "100111001010" => A <= "000000000000000000"; -- Line 157   Column 11   Coefficient 0.00000000
         when "100111001011" => A <= "000000000000000000"; -- Line 157   Column 12   Coefficient 0.00000000
         when "100111001100" => A <= "000000000000000000"; -- Line 157   Column 13   Coefficient 0.00000000
         when "100111001101" => A <= "000000000000000000"; -- Line 157   Column 14   Coefficient 0.00000000
         when "100111001110" => A <= "000000000000000000"; -- Line 157   Column 15   Coefficient 0.00000000
         when "100111001111" => A <= "000000000000000000"; -- Line 157   Column 16   Coefficient 0.00000000
         when "100111010000" => A <= "000000000000000000"; -- Line 158   Column 1   Coefficient 0.00000000
         when "100111010001" => A <= "000000000000000000"; -- Line 158   Column 2   Coefficient 0.00000000
         when "100111010010" => A <= "000000000000000000"; -- Line 158   Column 3   Coefficient 0.00000000
         when "100111010011" => A <= "000000000000000000"; -- Line 158   Column 4   Coefficient 0.00000000
         when "100111010100" => A <= "000000001111000010"; -- Line 158   Column 5   Coefficient 0.00366974
         when "100111010101" => A <= "111110000010011110"; -- Line 158   Column 6   Coefficient -0.03064728
         when "100111010110" => A <= "010011010010100110"; -- Line 158   Column 7   Coefficient 0.30141449
         when "100111010111" => A <= "111101100111001110"; -- Line 158   Column 8   Coefficient -0.03730011
         when "100111011000" => A <= "000000110010101110"; -- Line 158   Column 9   Coefficient 0.01238251
         when "100111011001" => A <= "000000000001111110"; -- Line 158   Column 10   Coefficient 0.00048065
         when "100111011010" => A <= "000000000000000000"; -- Line 158   Column 11   Coefficient 0.00000000
         when "100111011011" => A <= "000000000000000000"; -- Line 158   Column 12   Coefficient 0.00000000
         when "100111011100" => A <= "000000000000000000"; -- Line 158   Column 13   Coefficient 0.00000000
         when "100111011101" => A <= "000000000000000000"; -- Line 158   Column 14   Coefficient 0.00000000
         when "100111011110" => A <= "000000000000000000"; -- Line 158   Column 15   Coefficient 0.00000000
         when "100111011111" => A <= "000000000000000000"; -- Line 158   Column 16   Coefficient 0.00000000
         when "100111100000" => A <= "000000000000000000"; -- Line 159   Column 1   Coefficient 0.00000000
         when "100111100001" => A <= "000000000000000000"; -- Line 159   Column 2   Coefficient 0.00000000
         when "100111100010" => A <= "000000000000000000"; -- Line 159   Column 3   Coefficient 0.00000000
         when "100111100011" => A <= "000000000000000000"; -- Line 159   Column 4   Coefficient 0.00000000
         when "100111100100" => A <= "000000010000011000"; -- Line 159   Column 5   Coefficient 0.00399780
         when "100111100101" => A <= "111101101011101110"; -- Line 159   Column 6   Coefficient -0.03620148
         when "100111100110" => A <= "010010110100110100"; -- Line 159   Column 7   Coefficient 0.29414368
         when "100111100111" => A <= "111110100000101100"; -- Line 159   Column 8   Coefficient -0.02326965
         when "100111101000" => A <= "000000101101010111"; -- Line 159   Column 9   Coefficient 0.01107407
         when "100111101001" => A <= "000000000001000010"; -- Line 159   Column 10   Coefficient 0.00025177
         when "100111101010" => A <= "000000000000000000"; -- Line 159   Column 11   Coefficient 0.00000000
         when "100111101011" => A <= "000000000000000000"; -- Line 159   Column 12   Coefficient 0.00000000
         when "100111101100" => A <= "000000000000000000"; -- Line 159   Column 13   Coefficient 0.00000000
         when "100111101101" => A <= "000000000000000000"; -- Line 159   Column 14   Coefficient 0.00000000
         when "100111101110" => A <= "000000000000000000"; -- Line 159   Column 15   Coefficient 0.00000000
         when "100111101111" => A <= "000000000000000000"; -- Line 159   Column 16   Coefficient 0.00000000
         when "100111110000" => A <= "000000000000000000"; -- Line 160   Column 1   Coefficient 0.00000000
         when "100111110001" => A <= "000000000000000000"; -- Line 160   Column 2   Coefficient 0.00000000
         when "100111110010" => A <= "000000000000000000"; -- Line 160   Column 3   Coefficient 0.00000000
         when "100111110011" => A <= "000000000000000000"; -- Line 160   Column 4   Coefficient 0.00000000
         when "100111110100" => A <= "000000001111111100"; -- Line 160   Column 5   Coefficient 0.00389099
         when "100111110101" => A <= "111101100000101101"; -- Line 160   Column 6   Coefficient -0.03889084
         when "100111110110" => A <= "010010000001100011"; -- Line 160   Column 7   Coefficient 0.28162766
         when "100111110111" => A <= "111111101010001000"; -- Line 160   Column 8   Coefficient -0.00534058
         when "100111111000" => A <= "000000100010100100"; -- Line 160   Column 9   Coefficient 0.00843811
         when "100111111001" => A <= "000000000001001000"; -- Line 160   Column 10   Coefficient 0.00027466
         when "100111111010" => A <= "000000000000000000"; -- Line 160   Column 11   Coefficient 0.00000000
         when "100111111011" => A <= "000000000000000000"; -- Line 160   Column 12   Coefficient 0.00000000
         when "100111111100" => A <= "000000000000000000"; -- Line 160   Column 13   Coefficient 0.00000000
         when "100111111101" => A <= "000000000000000000"; -- Line 160   Column 14   Coefficient 0.00000000
         when "100111111110" => A <= "000000000000000000"; -- Line 160   Column 15   Coefficient 0.00000000
         when "100111111111" => A <= "000000000000000000"; -- Line 160   Column 16   Coefficient 0.00000000
         when "101000000000" => A <= "000000000000000000"; -- Line 161   Column 1   Coefficient 0.00000000
         when "101000000001" => A <= "000000000000000000"; -- Line 161   Column 2   Coefficient 0.00000000
         when "101000000010" => A <= "000000000000000000"; -- Line 161   Column 3   Coefficient 0.00000000
         when "101000000011" => A <= "000000000000000000"; -- Line 161   Column 4   Coefficient 0.00000000
         when "101000000100" => A <= "000000001101001100"; -- Line 161   Column 5   Coefficient 0.00321960
         when "101000000101" => A <= "111101100010001110"; -- Line 161   Column 6   Coefficient -0.03852081
         when "101000000110" => A <= "010000111010100101"; -- Line 161   Column 7   Coefficient 0.26430130
         when "101000000111" => A <= "000000111110100110"; -- Line 161   Column 8   Coefficient 0.01528168
         when "101000001000" => A <= "000000010110010000"; -- Line 161   Column 9   Coefficient 0.00543213
         when "101000001001" => A <= "000000000001001011"; -- Line 161   Column 10   Coefficient 0.00028610
         when "101000001010" => A <= "000000000000000000"; -- Line 161   Column 11   Coefficient 0.00000000
         when "101000001011" => A <= "000000000000000000"; -- Line 161   Column 12   Coefficient 0.00000000
         when "101000001100" => A <= "000000000000000000"; -- Line 161   Column 13   Coefficient 0.00000000
         when "101000001101" => A <= "000000000000000000"; -- Line 161   Column 14   Coefficient 0.00000000
         when "101000001110" => A <= "000000000000000000"; -- Line 161   Column 15   Coefficient 0.00000000
         when "101000001111" => A <= "000000000000000000"; -- Line 161   Column 16   Coefficient 0.00000000
         when "101000010000" => A <= "000000000000000000"; -- Line 162   Column 1   Coefficient 0.00000000
         when "101000010001" => A <= "000000000000000000"; -- Line 162   Column 2   Coefficient 0.00000000
         when "101000010010" => A <= "000000000000000000"; -- Line 162   Column 3   Coefficient 0.00000000
         when "101000010011" => A <= "000000000000000000"; -- Line 162   Column 4   Coefficient 0.00000000
         when "101000010100" => A <= "000000001010110110"; -- Line 162   Column 5   Coefficient 0.00264740
         when "101000010101" => A <= "111101100010101111"; -- Line 162   Column 6   Coefficient -0.03839493
         when "101000010110" => A <= "001111111010100001"; -- Line 162   Column 7   Coefficient 0.24866104
         when "101000010111" => A <= "000010000100001011"; -- Line 162   Column 8   Coefficient 0.03226852
         when "101000011000" => A <= "000000010100110111"; -- Line 162   Column 9   Coefficient 0.00509262
         when "101000011001" => A <= "111111111110110111"; -- Line 162   Column 10   Coefficient -0.00027847
         when "101000011010" => A <= "000000000000000000"; -- Line 162   Column 11   Coefficient 0.00000000
         when "101000011011" => A <= "000000000000000000"; -- Line 162   Column 12   Coefficient 0.00000000
         when "101000011100" => A <= "000000000000000000"; -- Line 162   Column 13   Coefficient 0.00000000
         when "101000011101" => A <= "000000000000000000"; -- Line 162   Column 14   Coefficient 0.00000000
         when "101000011110" => A <= "000000000000000000"; -- Line 162   Column 15   Coefficient 0.00000000
         when "101000011111" => A <= "000000000000000000"; -- Line 162   Column 16   Coefficient 0.00000000
         when "101000100000" => A <= "000000000000000000"; -- Line 163   Column 1   Coefficient 0.00000000
         when "101000100001" => A <= "000000000000000000"; -- Line 163   Column 2   Coefficient 0.00000000
         when "101000100010" => A <= "000000000000000000"; -- Line 163   Column 3   Coefficient 0.00000000
         when "101000100011" => A <= "000000000000000000"; -- Line 163   Column 4   Coefficient 0.00000000
         when "101000100100" => A <= "000000001000010011"; -- Line 163   Column 5   Coefficient 0.00202560
         when "101000100101" => A <= "111101100110110000"; -- Line 163   Column 6   Coefficient -0.03741455
         when "101000100110" => A <= "001110110101010100"; -- Line 163   Column 7   Coefficient 0.23176575
         when "101000100111" => A <= "000011001010010011"; -- Line 163   Column 8   Coefficient 0.04938889
         when "101000101000" => A <= "000000010100111001"; -- Line 163   Column 9   Coefficient 0.00510025
         when "101000101001" => A <= "111111111100011110"; -- Line 163   Column 10   Coefficient -0.00086212
         when "101000101010" => A <= "111111111111111111"; -- Line 163   Column 11   Coefficient -0.00000381
         when "101000101011" => A <= "000000000000000000"; -- Line 163   Column 12   Coefficient 0.00000000
         when "101000101100" => A <= "000000000000000000"; -- Line 163   Column 13   Coefficient 0.00000000
         when "101000101101" => A <= "000000000000000000"; -- Line 163   Column 14   Coefficient 0.00000000
         when "101000101110" => A <= "000000000000000000"; -- Line 163   Column 15   Coefficient 0.00000000
         when "101000101111" => A <= "000000000000000000"; -- Line 163   Column 16   Coefficient 0.00000000
         when "101000110000" => A <= "000000000000000000"; -- Line 164   Column 1   Coefficient 0.00000000
         when "101000110001" => A <= "000000000000000000"; -- Line 164   Column 2   Coefficient 0.00000000
         when "101000110010" => A <= "000000000000000000"; -- Line 164   Column 3   Coefficient 0.00000000
         when "101000110011" => A <= "000000000000000000"; -- Line 164   Column 4   Coefficient 0.00000000
         when "101000110100" => A <= "000000000011111000"; -- Line 164   Column 5   Coefficient 0.00094604
         when "101000110101" => A <= "111101110100001010"; -- Line 164   Column 6   Coefficient -0.03414154
         when "101000110110" => A <= "001101100011111111"; -- Line 164   Column 7   Coefficient 0.21191025
         when "101000110111" => A <= "000100010011001101"; -- Line 164   Column 8   Coefficient 0.06718826
         when "101000111000" => A <= "000000010111101010"; -- Line 164   Column 9   Coefficient 0.00577545
         when "101000111001" => A <= "111111111001000110"; -- Line 164   Column 10   Coefficient -0.00168610
         when "101000111010" => A <= "000000000000000011"; -- Line 164   Column 11   Coefficient 0.00001144
         when "101000111011" => A <= "000000000000000000"; -- Line 164   Column 12   Coefficient 0.00000000
         when "101000111100" => A <= "000000000000000000"; -- Line 164   Column 13   Coefficient 0.00000000
         when "101000111101" => A <= "000000000000000000"; -- Line 164   Column 14   Coefficient 0.00000000
         when "101000111110" => A <= "000000000000000000"; -- Line 164   Column 15   Coefficient 0.00000000
         when "101000111111" => A <= "000000000000000000"; -- Line 164   Column 16   Coefficient 0.00000000
         when "101001000000" => A <= "000000000000000000"; -- Line 165   Column 1   Coefficient 0.00000000
         when "101001000001" => A <= "000000000000000000"; -- Line 165   Column 2   Coefficient 0.00000000
         when "101001000010" => A <= "000000000000000000"; -- Line 165   Column 3   Coefficient 0.00000000
         when "101001000011" => A <= "000000000000000000"; -- Line 165   Column 4   Coefficient 0.00000000
         when "101001000100" => A <= "111111111111010011"; -- Line 165   Column 5   Coefficient -0.00017166
         when "101001000101" => A <= "111110000101010011"; -- Line 165   Column 6   Coefficient -0.02995682
         when "101001000110" => A <= "001100001011101000"; -- Line 165   Column 7   Coefficient 0.19033813
         when "101001000111" => A <= "000101100000010101"; -- Line 165   Column 8   Coefficient 0.08601761
         when "101001001000" => A <= "000000011000110111"; -- Line 165   Column 9   Coefficient 0.00606918
         when "101001001001" => A <= "111111110110011111"; -- Line 165   Column 10   Coefficient -0.00232315
         when "101001001010" => A <= "000000000000000110"; -- Line 165   Column 11   Coefficient 0.00002289
         when "101001001011" => A <= "000000000000000000"; -- Line 165   Column 12   Coefficient 0.00000000
         when "101001001100" => A <= "000000000000000000"; -- Line 165   Column 13   Coefficient 0.00000000
         when "101001001101" => A <= "000000000000000000"; -- Line 165   Column 14   Coefficient 0.00000000
         when "101001001110" => A <= "000000000000000000"; -- Line 165   Column 15   Coefficient 0.00000000
         when "101001001111" => A <= "000000000000000000"; -- Line 165   Column 16   Coefficient 0.00000000
         when "101001010000" => A <= "000000000000000000"; -- Line 166   Column 1   Coefficient 0.00000000
         when "101001010001" => A <= "000000000000000000"; -- Line 166   Column 2   Coefficient 0.00000000
         when "101001010010" => A <= "000000000000000000"; -- Line 166   Column 3   Coefficient 0.00000000
         when "101001010011" => A <= "000000000000000000"; -- Line 166   Column 4   Coefficient 0.00000000
         when "101001010100" => A <= "111111111110010010"; -- Line 166   Column 5   Coefficient -0.00041962
         when "101001010101" => A <= "111110010000110000"; -- Line 166   Column 6   Coefficient -0.02716064
         when "101001010110" => A <= "001010101100000111"; -- Line 166   Column 7   Coefficient 0.16701889
         when "101001010111" => A <= "000111000101010101"; -- Line 166   Column 8   Coefficient 0.11067581
         when "101001011000" => A <= "000000000100100100"; -- Line 166   Column 9   Coefficient 0.00111389
         when "101001011001" => A <= "111111111010111001"; -- Line 166   Column 10   Coefficient -0.00124741
         when "101001011010" => A <= "000000000000000100"; -- Line 166   Column 11   Coefficient 0.00001526
         when "101001011011" => A <= "000000000000000000"; -- Line 166   Column 12   Coefficient 0.00000000
         when "101001011100" => A <= "000000000000000000"; -- Line 166   Column 13   Coefficient 0.00000000
         when "101001011101" => A <= "000000000000000000"; -- Line 166   Column 14   Coefficient 0.00000000
         when "101001011110" => A <= "000000000000000000"; -- Line 166   Column 15   Coefficient 0.00000000
         when "101001011111" => A <= "000000000000000000"; -- Line 166   Column 16   Coefficient 0.00000000
         when "101001100000" => A <= "000000000000000000"; -- Line 167   Column 1   Coefficient 0.00000000
         when "101001100001" => A <= "000000000000000000"; -- Line 167   Column 2   Coefficient 0.00000000
         when "101001100010" => A <= "000000000000000000"; -- Line 167   Column 3   Coefficient 0.00000000
         when "101001100011" => A <= "000000000000000000"; -- Line 167   Column 4   Coefficient 0.00000000
         when "101001100100" => A <= "111111111110100110"; -- Line 167   Column 5   Coefficient -0.00034332
         when "101001100101" => A <= "111110011011111010"; -- Line 167   Column 6   Coefficient -0.02443695
         when "101001100110" => A <= "001001000110101001"; -- Line 167   Column 7   Coefficient 0.14224625
         when "101001100111" => A <= "001000110101000000"; -- Line 167   Column 8   Coefficient 0.13793945
         when "101001101000" => A <= "111111100111100010"; -- Line 167   Column 9   Coefficient -0.00597382
         when "101001101001" => A <= "000000000010010011"; -- Line 167   Column 10   Coefficient 0.00056076
         when "101001101010" => A <= "000000000000000011"; -- Line 167   Column 11   Coefficient 0.00001144
         when "101001101011" => A <= "000000000000000000"; -- Line 167   Column 12   Coefficient 0.00000000
         when "101001101100" => A <= "000000000000000000"; -- Line 167   Column 13   Coefficient 0.00000000
         when "101001101101" => A <= "000000000000000000"; -- Line 167   Column 14   Coefficient 0.00000000
         when "101001101110" => A <= "000000000000000000"; -- Line 167   Column 15   Coefficient 0.00000000
         when "101001101111" => A <= "000000000000000000"; -- Line 167   Column 16   Coefficient 0.00000000
         when "101001110000" => A <= "000000000000000000"; -- Line 168   Column 1   Coefficient 0.00000000
         when "101001110001" => A <= "000000000000000000"; -- Line 168   Column 2   Coefficient 0.00000000
         when "101001110010" => A <= "000000000000000000"; -- Line 168   Column 3   Coefficient 0.00000000
         when "101001110011" => A <= "000000000000000000"; -- Line 168   Column 4   Coefficient 0.00000000
         when "101001110100" => A <= "111111111111001011"; -- Line 168   Column 5   Coefficient -0.00020218
         when "101001110101" => A <= "111110100110010011"; -- Line 168   Column 6   Coefficient -0.02190018
         when "101001110110" => A <= "000111100110110001"; -- Line 168   Column 7   Coefficient 0.11883926
         when "101001110111" => A <= "001010011001111000"; -- Line 168   Column 8   Coefficient 0.16256714
         when "101001111000" => A <= "111111010000101110"; -- Line 168   Column 9   Coefficient -0.01154327
         when "101001111001" => A <= "000000001001011000"; -- Line 168   Column 10   Coefficient 0.00228882
         when "101001111010" => A <= "111111111111110100"; -- Line 168   Column 11   Coefficient -0.00004578
         when "101001111011" => A <= "000000000000000000"; -- Line 168   Column 12   Coefficient 0.00000000
         when "101001111100" => A <= "000000000000000000"; -- Line 168   Column 13   Coefficient 0.00000000
         when "101001111101" => A <= "000000000000000000"; -- Line 168   Column 14   Coefficient 0.00000000
         when "101001111110" => A <= "000000000000000000"; -- Line 168   Column 15   Coefficient 0.00000000
         when "101001111111" => A <= "000000000000000000"; -- Line 168   Column 16   Coefficient 0.00000000
         when "101010000000" => A <= "000000000000000000"; -- Line 169   Column 1   Coefficient 0.00000000
         when "101010000001" => A <= "000000000000000000"; -- Line 169   Column 2   Coefficient 0.00000000
         when "101010000010" => A <= "000000000000000000"; -- Line 169   Column 3   Coefficient 0.00000000
         when "101010000011" => A <= "000000000000000000"; -- Line 169   Column 4   Coefficient 0.00000000
         when "101010000100" => A <= "000000000000000011"; -- Line 169   Column 5   Coefficient 0.00001144
         when "101010000101" => A <= "111110110001100001"; -- Line 169   Column 6   Coefficient -0.01916122
         when "101010000110" => A <= "000110000101110011"; -- Line 169   Column 7   Coefficient 0.09516525
         when "101010000111" => A <= "001011111101111010"; -- Line 169   Column 8   Coefficient 0.18698883
         when "101010001000" => A <= "111110111010000001"; -- Line 169   Column 9   Coefficient -0.01708603
         when "101010001001" => A <= "000000010001001000"; -- Line 169   Column 10   Coefficient 0.00418091
         when "101010001010" => A <= "111111111111100110"; -- Line 169   Column 11   Coefficient -0.00009918
         when "101010001011" => A <= "000000000000000000"; -- Line 169   Column 12   Coefficient 0.00000000
         when "101010001100" => A <= "000000000000000000"; -- Line 169   Column 13   Coefficient 0.00000000
         when "101010001101" => A <= "000000000000000000"; -- Line 169   Column 14   Coefficient 0.00000000
         when "101010001110" => A <= "000000000000000000"; -- Line 169   Column 15   Coefficient 0.00000000
         when "101010001111" => A <= "000000000000000000"; -- Line 169   Column 16   Coefficient 0.00000000
         when "101010010000" => A <= "000000000000000000"; -- Line 170   Column 1   Coefficient 0.00000000
         when "101010010001" => A <= "000000000000000000"; -- Line 170   Column 2   Coefficient 0.00000000
         when "101010010010" => A <= "000000000000000000"; -- Line 170   Column 3   Coefficient 0.00000000
         when "101010010011" => A <= "000000000000000000"; -- Line 170   Column 4   Coefficient 0.00000000
         when "101010010100" => A <= "000000000000001001"; -- Line 170   Column 5   Coefficient 0.00003433
         when "101010010101" => A <= "111111000100111001"; -- Line 170   Column 6   Coefficient -0.01443100
         when "101010010110" => A <= "000100010010000101"; -- Line 170   Column 7   Coefficient 0.06691360
         when "101010010111" => A <= "001101110100101001"; -- Line 170   Column 8   Coefficient 0.21597672
         when "101010011000" => A <= "111110011010010101"; -- Line 170   Column 9   Coefficient -0.02482224
         when "101010011001" => A <= "000000011001110100"; -- Line 170   Column 10   Coefficient 0.00630188
         when "101010011010" => A <= "000000000000000111"; -- Line 170   Column 11   Coefficient 0.00002670
         when "101010011011" => A <= "000000000000000000"; -- Line 170   Column 12   Coefficient 0.00000000
         when "101010011100" => A <= "000000000000000000"; -- Line 170   Column 13   Coefficient 0.00000000
         when "101010011101" => A <= "000000000000000000"; -- Line 170   Column 14   Coefficient 0.00000000
         when "101010011110" => A <= "000000000000000000"; -- Line 170   Column 15   Coefficient 0.00000000
         when "101010011111" => A <= "000000000000000000"; -- Line 170   Column 16   Coefficient 0.00000000
         when "101010100000" => A <= "000000000000000000"; -- Line 171   Column 1   Coefficient 0.00000000
         when "101010100001" => A <= "000000000000000000"; -- Line 171   Column 2   Coefficient 0.00000000
         when "101010100010" => A <= "000000000000000000"; -- Line 171   Column 3   Coefficient 0.00000000
         when "101010100011" => A <= "000000000000000000"; -- Line 171   Column 4   Coefficient 0.00000000
         when "101010100100" => A <= "000000000000000000"; -- Line 171   Column 5   Coefficient 0.00000000
         when "101010100101" => A <= "111111011001111001"; -- Line 171   Column 6   Coefficient -0.00930405
         when "101010100110" => A <= "000010011110111100"; -- Line 171   Column 7   Coefficient 0.03880310
         when "101010100111" => A <= "001111100101110011"; -- Line 171   Column 8   Coefficient 0.24360275
         when "101010101000" => A <= "111101111110110001"; -- Line 171   Column 9   Coefficient -0.03155136
         when "101010101001" => A <= "000000100001110011"; -- Line 171   Column 10   Coefficient 0.00825119
         when "101010101010" => A <= "000000000000110011"; -- Line 171   Column 11   Coefficient 0.00019455
         when "101010101011" => A <= "000000000000000000"; -- Line 171   Column 12   Coefficient 0.00000000
         when "101010101100" => A <= "000000000000000000"; -- Line 171   Column 13   Coefficient 0.00000000
         when "101010101101" => A <= "000000000000000000"; -- Line 171   Column 14   Coefficient 0.00000000
         when "101010101110" => A <= "000000000000000000"; -- Line 171   Column 15   Coefficient 0.00000000
         when "101010101111" => A <= "000000000000000000"; -- Line 171   Column 16   Coefficient 0.00000000
         when "101010110000" => A <= "000000000000000000"; -- Line 172   Column 1   Coefficient 0.00000000
         when "101010110001" => A <= "000000000000000000"; -- Line 172   Column 2   Coefficient 0.00000000
         when "101010110010" => A <= "000000000000000000"; -- Line 172   Column 3   Coefficient 0.00000000
         when "101010110011" => A <= "000000000000000000"; -- Line 172   Column 4   Coefficient 0.00000000
         when "101010110100" => A <= "000000000000000000"; -- Line 172   Column 5   Coefficient 0.00000000
         when "101010110101" => A <= "111111110001010101"; -- Line 172   Column 6   Coefficient -0.00358200
         when "101010110110" => A <= "000000100101011001"; -- Line 172   Column 7   Coefficient 0.00912857
         when "101010110111" => A <= "010001011110001011"; -- Line 172   Column 8   Coefficient 0.27299118
         when "101010111000" => A <= "111101011101101101"; -- Line 172   Column 9   Coefficient -0.03962326
         when "101010111001" => A <= "000000101011110101"; -- Line 172   Column 10   Coefficient 0.01070023
         when "101010111010" => A <= "000000000001100101"; -- Line 172   Column 11   Coefficient 0.00038528
         when "101010111011" => A <= "000000000000000000"; -- Line 172   Column 12   Coefficient 0.00000000
         when "101010111100" => A <= "000000000000000000"; -- Line 172   Column 13   Coefficient 0.00000000
         when "101010111101" => A <= "000000000000000000"; -- Line 172   Column 14   Coefficient 0.00000000
         when "101010111110" => A <= "000000000000000000"; -- Line 172   Column 15   Coefficient 0.00000000
         when "101010111111" => A <= "000000000000000000"; -- Line 172   Column 16   Coefficient 0.00000000
         when "101011000000" => A <= "000000000000000000"; -- Line 173   Column 1   Coefficient 0.00000000
         when "101011000001" => A <= "000000000000000000"; -- Line 173   Column 2   Coefficient 0.00000000
         when "101011000010" => A <= "000000000000000000"; -- Line 173   Column 3   Coefficient 0.00000000
         when "101011000011" => A <= "000000000000000000"; -- Line 173   Column 4   Coefficient 0.00000000
         when "101011000100" => A <= "000000000000000000"; -- Line 173   Column 5   Coefficient 0.00000000
         when "101011000101" => A <= "000000000111011010"; -- Line 173   Column 6   Coefficient 0.00180817
         when "101011000110" => A <= "111110110101100100"; -- Line 173   Column 7   Coefficient -0.01817322
         when "101011000111" => A <= "010011000101100111"; -- Line 173   Column 8   Coefficient 0.29824448
         when "101011001000" => A <= "111101000110110001"; -- Line 173   Column 9   Coefficient -0.04522324
         when "101011001001" => A <= "000000110100010110"; -- Line 173   Column 10   Coefficient 0.01277924
         when "101011001010" => A <= "000000000010010101"; -- Line 173   Column 11   Coefficient 0.00056839
         when "101011001011" => A <= "000000000000000000"; -- Line 173   Column 12   Coefficient 0.00000000
         when "101011001100" => A <= "000000000000000000"; -- Line 173   Column 13   Coefficient 0.00000000
         when "101011001101" => A <= "000000000000000000"; -- Line 173   Column 14   Coefficient 0.00000000
         when "101011001110" => A <= "000000000000000000"; -- Line 173   Column 15   Coefficient 0.00000000
         when "101011001111" => A <= "000000000000000000"; -- Line 173   Column 16   Coefficient 0.00000000
         when "101011010000" => A <= "000000000000000000"; -- Line 174   Column 1   Coefficient 0.00000000
         when "101011010001" => A <= "000000000000000000"; -- Line 174   Column 2   Coefficient 0.00000000
         when "101011010010" => A <= "000000000000000000"; -- Line 174   Column 3   Coefficient 0.00000000
         when "101011010011" => A <= "000000000000000000"; -- Line 174   Column 4   Coefficient 0.00000000
         when "101011010100" => A <= "000000000000000000"; -- Line 174   Column 5   Coefficient 0.00000000
         when "101011010101" => A <= "000000001111000010"; -- Line 174   Column 6   Coefficient 0.00366974
         when "101011010110" => A <= "111110000010011110"; -- Line 174   Column 7   Coefficient -0.03064728
         when "101011010111" => A <= "010011010010100110"; -- Line 174   Column 8   Coefficient 0.30141449
         when "101011011000" => A <= "111101100111001110"; -- Line 174   Column 9   Coefficient -0.03730011
         when "101011011001" => A <= "000000110010101110"; -- Line 174   Column 10   Coefficient 0.01238251
         when "101011011010" => A <= "000000000001111110"; -- Line 174   Column 11   Coefficient 0.00048065
         when "101011011011" => A <= "000000000000000000"; -- Line 174   Column 12   Coefficient 0.00000000
         when "101011011100" => A <= "000000000000000000"; -- Line 174   Column 13   Coefficient 0.00000000
         when "101011011101" => A <= "000000000000000000"; -- Line 174   Column 14   Coefficient 0.00000000
         when "101011011110" => A <= "000000000000000000"; -- Line 174   Column 15   Coefficient 0.00000000
         when "101011011111" => A <= "000000000000000000"; -- Line 174   Column 16   Coefficient 0.00000000
         when "101011100000" => A <= "000000000000000000"; -- Line 175   Column 1   Coefficient 0.00000000
         when "101011100001" => A <= "000000000000000000"; -- Line 175   Column 2   Coefficient 0.00000000
         when "101011100010" => A <= "000000000000000000"; -- Line 175   Column 3   Coefficient 0.00000000
         when "101011100011" => A <= "000000000000000000"; -- Line 175   Column 4   Coefficient 0.00000000
         when "101011100100" => A <= "000000000000000000"; -- Line 175   Column 5   Coefficient 0.00000000
         when "101011100101" => A <= "000000010000011000"; -- Line 175   Column 6   Coefficient 0.00399780
         when "101011100110" => A <= "111101101011101110"; -- Line 175   Column 7   Coefficient -0.03620148
         when "101011100111" => A <= "010010110100110100"; -- Line 175   Column 8   Coefficient 0.29414368
         when "101011101000" => A <= "111110100000101100"; -- Line 175   Column 9   Coefficient -0.02326965
         when "101011101001" => A <= "000000101101010111"; -- Line 175   Column 10   Coefficient 0.01107407
         when "101011101010" => A <= "000000000001000010"; -- Line 175   Column 11   Coefficient 0.00025177
         when "101011101011" => A <= "000000000000000000"; -- Line 175   Column 12   Coefficient 0.00000000
         when "101011101100" => A <= "000000000000000000"; -- Line 175   Column 13   Coefficient 0.00000000
         when "101011101101" => A <= "000000000000000000"; -- Line 175   Column 14   Coefficient 0.00000000
         when "101011101110" => A <= "000000000000000000"; -- Line 175   Column 15   Coefficient 0.00000000
         when "101011101111" => A <= "000000000000000000"; -- Line 175   Column 16   Coefficient 0.00000000
         when "101011110000" => A <= "000000000000000000"; -- Line 176   Column 1   Coefficient 0.00000000
         when "101011110001" => A <= "000000000000000000"; -- Line 176   Column 2   Coefficient 0.00000000
         when "101011110010" => A <= "000000000000000000"; -- Line 176   Column 3   Coefficient 0.00000000
         when "101011110011" => A <= "000000000000000000"; -- Line 176   Column 4   Coefficient 0.00000000
         when "101011110100" => A <= "000000000000000000"; -- Line 176   Column 5   Coefficient 0.00000000
         when "101011110101" => A <= "000000001111111100"; -- Line 176   Column 6   Coefficient 0.00389099
         when "101011110110" => A <= "111101100000101101"; -- Line 176   Column 7   Coefficient -0.03889084
         when "101011110111" => A <= "010010000001100011"; -- Line 176   Column 8   Coefficient 0.28162766
         when "101011111000" => A <= "111111101010001000"; -- Line 176   Column 9   Coefficient -0.00534058
         when "101011111001" => A <= "000000100010100100"; -- Line 176   Column 10   Coefficient 0.00843811
         when "101011111010" => A <= "000000000001001000"; -- Line 176   Column 11   Coefficient 0.00027466
         when "101011111011" => A <= "000000000000000000"; -- Line 176   Column 12   Coefficient 0.00000000
         when "101011111100" => A <= "000000000000000000"; -- Line 176   Column 13   Coefficient 0.00000000
         when "101011111101" => A <= "000000000000000000"; -- Line 176   Column 14   Coefficient 0.00000000
         when "101011111110" => A <= "000000000000000000"; -- Line 176   Column 15   Coefficient 0.00000000
         when "101011111111" => A <= "000000000000000000"; -- Line 176   Column 16   Coefficient 0.00000000
         when "101100000000" => A <= "000000000000000000"; -- Line 177   Column 1   Coefficient 0.00000000
         when "101100000001" => A <= "000000000000000000"; -- Line 177   Column 2   Coefficient 0.00000000
         when "101100000010" => A <= "000000000000000000"; -- Line 177   Column 3   Coefficient 0.00000000
         when "101100000011" => A <= "000000000000000000"; -- Line 177   Column 4   Coefficient 0.00000000
         when "101100000100" => A <= "000000000000000000"; -- Line 177   Column 5   Coefficient 0.00000000
         when "101100000101" => A <= "000000001101001100"; -- Line 177   Column 6   Coefficient 0.00321960
         when "101100000110" => A <= "111101100010001110"; -- Line 177   Column 7   Coefficient -0.03852081
         when "101100000111" => A <= "010000111010100101"; -- Line 177   Column 8   Coefficient 0.26430130
         when "101100001000" => A <= "000000111110100110"; -- Line 177   Column 9   Coefficient 0.01528168
         when "101100001001" => A <= "000000010110010000"; -- Line 177   Column 10   Coefficient 0.00543213
         when "101100001010" => A <= "000000000001001011"; -- Line 177   Column 11   Coefficient 0.00028610
         when "101100001011" => A <= "000000000000000000"; -- Line 177   Column 12   Coefficient 0.00000000
         when "101100001100" => A <= "000000000000000000"; -- Line 177   Column 13   Coefficient 0.00000000
         when "101100001101" => A <= "000000000000000000"; -- Line 177   Column 14   Coefficient 0.00000000
         when "101100001110" => A <= "000000000000000000"; -- Line 177   Column 15   Coefficient 0.00000000
         when "101100001111" => A <= "000000000000000000"; -- Line 177   Column 16   Coefficient 0.00000000
         when "101100010000" => A <= "000000000000000000"; -- Line 178   Column 1   Coefficient 0.00000000
         when "101100010001" => A <= "000000000000000000"; -- Line 178   Column 2   Coefficient 0.00000000
         when "101100010010" => A <= "000000000000000000"; -- Line 178   Column 3   Coefficient 0.00000000
         when "101100010011" => A <= "000000000000000000"; -- Line 178   Column 4   Coefficient 0.00000000
         when "101100010100" => A <= "000000000000000000"; -- Line 178   Column 5   Coefficient 0.00000000
         when "101100010101" => A <= "000000001010110110"; -- Line 178   Column 6   Coefficient 0.00264740
         when "101100010110" => A <= "111101100010101111"; -- Line 178   Column 7   Coefficient -0.03839493
         when "101100010111" => A <= "001111111010100001"; -- Line 178   Column 8   Coefficient 0.24866104
         when "101100011000" => A <= "000010000100001011"; -- Line 178   Column 9   Coefficient 0.03226852
         when "101100011001" => A <= "000000010100110111"; -- Line 178   Column 10   Coefficient 0.00509262
         when "101100011010" => A <= "111111111110110111"; -- Line 178   Column 11   Coefficient -0.00027847
         when "101100011011" => A <= "000000000000000000"; -- Line 178   Column 12   Coefficient 0.00000000
         when "101100011100" => A <= "000000000000000000"; -- Line 178   Column 13   Coefficient 0.00000000
         when "101100011101" => A <= "000000000000000000"; -- Line 178   Column 14   Coefficient 0.00000000
         when "101100011110" => A <= "000000000000000000"; -- Line 178   Column 15   Coefficient 0.00000000
         when "101100011111" => A <= "000000000000000000"; -- Line 178   Column 16   Coefficient 0.00000000
         when "101100100000" => A <= "000000000000000000"; -- Line 179   Column 1   Coefficient 0.00000000
         when "101100100001" => A <= "000000000000000000"; -- Line 179   Column 2   Coefficient 0.00000000
         when "101100100010" => A <= "000000000000000000"; -- Line 179   Column 3   Coefficient 0.00000000
         when "101100100011" => A <= "000000000000000000"; -- Line 179   Column 4   Coefficient 0.00000000
         when "101100100100" => A <= "000000000000000000"; -- Line 179   Column 5   Coefficient 0.00000000
         when "101100100101" => A <= "000000001000010011"; -- Line 179   Column 6   Coefficient 0.00202560
         when "101100100110" => A <= "111101100110110000"; -- Line 179   Column 7   Coefficient -0.03741455
         when "101100100111" => A <= "001110110101010100"; -- Line 179   Column 8   Coefficient 0.23176575
         when "101100101000" => A <= "000011001010010011"; -- Line 179   Column 9   Coefficient 0.04938889
         when "101100101001" => A <= "000000010100111001"; -- Line 179   Column 10   Coefficient 0.00510025
         when "101100101010" => A <= "111111111100011110"; -- Line 179   Column 11   Coefficient -0.00086212
         when "101100101011" => A <= "111111111111111111"; -- Line 179   Column 12   Coefficient -0.00000381
         when "101100101100" => A <= "000000000000000000"; -- Line 179   Column 13   Coefficient 0.00000000
         when "101100101101" => A <= "000000000000000000"; -- Line 179   Column 14   Coefficient 0.00000000
         when "101100101110" => A <= "000000000000000000"; -- Line 179   Column 15   Coefficient 0.00000000
         when "101100101111" => A <= "000000000000000000"; -- Line 179   Column 16   Coefficient 0.00000000
         when "101100110000" => A <= "000000000000000000"; -- Line 180   Column 1   Coefficient 0.00000000
         when "101100110001" => A <= "000000000000000000"; -- Line 180   Column 2   Coefficient 0.00000000
         when "101100110010" => A <= "000000000000000000"; -- Line 180   Column 3   Coefficient 0.00000000
         when "101100110011" => A <= "000000000000000000"; -- Line 180   Column 4   Coefficient 0.00000000
         when "101100110100" => A <= "000000000000000000"; -- Line 180   Column 5   Coefficient 0.00000000
         when "101100110101" => A <= "000000000011111000"; -- Line 180   Column 6   Coefficient 0.00094604
         when "101100110110" => A <= "111101110100001010"; -- Line 180   Column 7   Coefficient -0.03414154
         when "101100110111" => A <= "001101100011111111"; -- Line 180   Column 8   Coefficient 0.21191025
         when "101100111000" => A <= "000100010011001101"; -- Line 180   Column 9   Coefficient 0.06718826
         when "101100111001" => A <= "000000010111101010"; -- Line 180   Column 10   Coefficient 0.00577545
         when "101100111010" => A <= "111111111001000110"; -- Line 180   Column 11   Coefficient -0.00168610
         when "101100111011" => A <= "000000000000000011"; -- Line 180   Column 12   Coefficient 0.00001144
         when "101100111100" => A <= "000000000000000000"; -- Line 180   Column 13   Coefficient 0.00000000
         when "101100111101" => A <= "000000000000000000"; -- Line 180   Column 14   Coefficient 0.00000000
         when "101100111110" => A <= "000000000000000000"; -- Line 180   Column 15   Coefficient 0.00000000
         when "101100111111" => A <= "000000000000000000"; -- Line 180   Column 16   Coefficient 0.00000000
         when "101101000000" => A <= "000000000000000000"; -- Line 181   Column 1   Coefficient 0.00000000
         when "101101000001" => A <= "000000000000000000"; -- Line 181   Column 2   Coefficient 0.00000000
         when "101101000010" => A <= "000000000000000000"; -- Line 181   Column 3   Coefficient 0.00000000
         when "101101000011" => A <= "000000000000000000"; -- Line 181   Column 4   Coefficient 0.00000000
         when "101101000100" => A <= "000000000000000000"; -- Line 181   Column 5   Coefficient 0.00000000
         when "101101000101" => A <= "111111111111010011"; -- Line 181   Column 6   Coefficient -0.00017166
         when "101101000110" => A <= "111110000101010011"; -- Line 181   Column 7   Coefficient -0.02995682
         when "101101000111" => A <= "001100001011101000"; -- Line 181   Column 8   Coefficient 0.19033813
         when "101101001000" => A <= "000101100000010101"; -- Line 181   Column 9   Coefficient 0.08601761
         when "101101001001" => A <= "000000011000110111"; -- Line 181   Column 10   Coefficient 0.00606918
         when "101101001010" => A <= "111111110110011111"; -- Line 181   Column 11   Coefficient -0.00232315
         when "101101001011" => A <= "000000000000000110"; -- Line 181   Column 12   Coefficient 0.00002289
         when "101101001100" => A <= "000000000000000000"; -- Line 181   Column 13   Coefficient 0.00000000
         when "101101001101" => A <= "000000000000000000"; -- Line 181   Column 14   Coefficient 0.00000000
         when "101101001110" => A <= "000000000000000000"; -- Line 181   Column 15   Coefficient 0.00000000
         when "101101001111" => A <= "000000000000000000"; -- Line 181   Column 16   Coefficient 0.00000000
         when "101101010000" => A <= "000000000000000000"; -- Line 182   Column 1   Coefficient 0.00000000
         when "101101010001" => A <= "000000000000000000"; -- Line 182   Column 2   Coefficient 0.00000000
         when "101101010010" => A <= "000000000000000000"; -- Line 182   Column 3   Coefficient 0.00000000
         when "101101010011" => A <= "000000000000000000"; -- Line 182   Column 4   Coefficient 0.00000000
         when "101101010100" => A <= "000000000000000000"; -- Line 182   Column 5   Coefficient 0.00000000
         when "101101010101" => A <= "111111111110010010"; -- Line 182   Column 6   Coefficient -0.00041962
         when "101101010110" => A <= "111110010000110000"; -- Line 182   Column 7   Coefficient -0.02716064
         when "101101010111" => A <= "001010101100000111"; -- Line 182   Column 8   Coefficient 0.16701889
         when "101101011000" => A <= "000111000101010101"; -- Line 182   Column 9   Coefficient 0.11067581
         when "101101011001" => A <= "000000000100100100"; -- Line 182   Column 10   Coefficient 0.00111389
         when "101101011010" => A <= "111111111010111001"; -- Line 182   Column 11   Coefficient -0.00124741
         when "101101011011" => A <= "000000000000000100"; -- Line 182   Column 12   Coefficient 0.00001526
         when "101101011100" => A <= "000000000000000000"; -- Line 182   Column 13   Coefficient 0.00000000
         when "101101011101" => A <= "000000000000000000"; -- Line 182   Column 14   Coefficient 0.00000000
         when "101101011110" => A <= "000000000000000000"; -- Line 182   Column 15   Coefficient 0.00000000
         when "101101011111" => A <= "000000000000000000"; -- Line 182   Column 16   Coefficient 0.00000000
         when "101101100000" => A <= "000000000000000000"; -- Line 183   Column 1   Coefficient 0.00000000
         when "101101100001" => A <= "000000000000000000"; -- Line 183   Column 2   Coefficient 0.00000000
         when "101101100010" => A <= "000000000000000000"; -- Line 183   Column 3   Coefficient 0.00000000
         when "101101100011" => A <= "000000000000000000"; -- Line 183   Column 4   Coefficient 0.00000000
         when "101101100100" => A <= "000000000000000000"; -- Line 183   Column 5   Coefficient 0.00000000
         when "101101100101" => A <= "111111111110100110"; -- Line 183   Column 6   Coefficient -0.00034332
         when "101101100110" => A <= "111110011011111010"; -- Line 183   Column 7   Coefficient -0.02443695
         when "101101100111" => A <= "001001000110101001"; -- Line 183   Column 8   Coefficient 0.14224625
         when "101101101000" => A <= "001000110101000000"; -- Line 183   Column 9   Coefficient 0.13793945
         when "101101101001" => A <= "111111100111100010"; -- Line 183   Column 10   Coefficient -0.00597382
         when "101101101010" => A <= "000000000010010011"; -- Line 183   Column 11   Coefficient 0.00056076
         when "101101101011" => A <= "000000000000000011"; -- Line 183   Column 12   Coefficient 0.00001144
         when "101101101100" => A <= "000000000000000000"; -- Line 183   Column 13   Coefficient 0.00000000
         when "101101101101" => A <= "000000000000000000"; -- Line 183   Column 14   Coefficient 0.00000000
         when "101101101110" => A <= "000000000000000000"; -- Line 183   Column 15   Coefficient 0.00000000
         when "101101101111" => A <= "000000000000000000"; -- Line 183   Column 16   Coefficient 0.00000000
         when "101101110000" => A <= "000000000000000000"; -- Line 184   Column 1   Coefficient 0.00000000
         when "101101110001" => A <= "000000000000000000"; -- Line 184   Column 2   Coefficient 0.00000000
         when "101101110010" => A <= "000000000000000000"; -- Line 184   Column 3   Coefficient 0.00000000
         when "101101110011" => A <= "000000000000000000"; -- Line 184   Column 4   Coefficient 0.00000000
         when "101101110100" => A <= "000000000000000000"; -- Line 184   Column 5   Coefficient 0.00000000
         when "101101110101" => A <= "111111111111001011"; -- Line 184   Column 6   Coefficient -0.00020218
         when "101101110110" => A <= "111110100110010011"; -- Line 184   Column 7   Coefficient -0.02190018
         when "101101110111" => A <= "000111100110110001"; -- Line 184   Column 8   Coefficient 0.11883926
         when "101101111000" => A <= "001010011001111000"; -- Line 184   Column 9   Coefficient 0.16256714
         when "101101111001" => A <= "111111010000101110"; -- Line 184   Column 10   Coefficient -0.01154327
         when "101101111010" => A <= "000000001001011000"; -- Line 184   Column 11   Coefficient 0.00228882
         when "101101111011" => A <= "111111111111110100"; -- Line 184   Column 12   Coefficient -0.00004578
         when "101101111100" => A <= "000000000000000000"; -- Line 184   Column 13   Coefficient 0.00000000
         when "101101111101" => A <= "000000000000000000"; -- Line 184   Column 14   Coefficient 0.00000000
         when "101101111110" => A <= "000000000000000000"; -- Line 184   Column 15   Coefficient 0.00000000
         when "101101111111" => A <= "000000000000000000"; -- Line 184   Column 16   Coefficient 0.00000000
         when "101110000000" => A <= "000000000000000000"; -- Line 185   Column 1   Coefficient 0.00000000
         when "101110000001" => A <= "000000000000000000"; -- Line 185   Column 2   Coefficient 0.00000000
         when "101110000010" => A <= "000000000000000000"; -- Line 185   Column 3   Coefficient 0.00000000
         when "101110000011" => A <= "000000000000000000"; -- Line 185   Column 4   Coefficient 0.00000000
         when "101110000100" => A <= "000000000000000000"; -- Line 185   Column 5   Coefficient 0.00000000
         when "101110000101" => A <= "000000000000000011"; -- Line 185   Column 6   Coefficient 0.00001144
         when "101110000110" => A <= "111110110001100001"; -- Line 185   Column 7   Coefficient -0.01916122
         when "101110000111" => A <= "000110000101110011"; -- Line 185   Column 8   Coefficient 0.09516525
         when "101110001000" => A <= "001011111101111010"; -- Line 185   Column 9   Coefficient 0.18698883
         when "101110001001" => A <= "111110111010000001"; -- Line 185   Column 10   Coefficient -0.01708603
         when "101110001010" => A <= "000000010001001000"; -- Line 185   Column 11   Coefficient 0.00418091
         when "101110001011" => A <= "111111111111100110"; -- Line 185   Column 12   Coefficient -0.00009918
         when "101110001100" => A <= "000000000000000000"; -- Line 185   Column 13   Coefficient 0.00000000
         when "101110001101" => A <= "000000000000000000"; -- Line 185   Column 14   Coefficient 0.00000000
         when "101110001110" => A <= "000000000000000000"; -- Line 185   Column 15   Coefficient 0.00000000
         when "101110001111" => A <= "000000000000000000"; -- Line 185   Column 16   Coefficient 0.00000000
         when "101110010000" => A <= "000000000000000000"; -- Line 186   Column 1   Coefficient 0.00000000
         when "101110010001" => A <= "000000000000000000"; -- Line 186   Column 2   Coefficient 0.00000000
         when "101110010010" => A <= "000000000000000000"; -- Line 186   Column 3   Coefficient 0.00000000
         when "101110010011" => A <= "000000000000000000"; -- Line 186   Column 4   Coefficient 0.00000000
         when "101110010100" => A <= "000000000000000000"; -- Line 186   Column 5   Coefficient 0.00000000
         when "101110010101" => A <= "000000000000001001"; -- Line 186   Column 6   Coefficient 0.00003433
         when "101110010110" => A <= "111111000100111001"; -- Line 186   Column 7   Coefficient -0.01443100
         when "101110010111" => A <= "000100010010000101"; -- Line 186   Column 8   Coefficient 0.06691360
         when "101110011000" => A <= "001101110100101001"; -- Line 186   Column 9   Coefficient 0.21597672
         when "101110011001" => A <= "111110011010010101"; -- Line 186   Column 10   Coefficient -0.02482224
         when "101110011010" => A <= "000000011001110100"; -- Line 186   Column 11   Coefficient 0.00630188
         when "101110011011" => A <= "000000000000000111"; -- Line 186   Column 12   Coefficient 0.00002670
         when "101110011100" => A <= "000000000000000000"; -- Line 186   Column 13   Coefficient 0.00000000
         when "101110011101" => A <= "000000000000000000"; -- Line 186   Column 14   Coefficient 0.00000000
         when "101110011110" => A <= "000000000000000000"; -- Line 186   Column 15   Coefficient 0.00000000
         when "101110011111" => A <= "000000000000000000"; -- Line 186   Column 16   Coefficient 0.00000000
         when "101110100000" => A <= "000000000000000000"; -- Line 187   Column 1   Coefficient 0.00000000
         when "101110100001" => A <= "000000000000000000"; -- Line 187   Column 2   Coefficient 0.00000000
         when "101110100010" => A <= "000000000000000000"; -- Line 187   Column 3   Coefficient 0.00000000
         when "101110100011" => A <= "000000000000000000"; -- Line 187   Column 4   Coefficient 0.00000000
         when "101110100100" => A <= "000000000000000000"; -- Line 187   Column 5   Coefficient 0.00000000
         when "101110100101" => A <= "000000000000000000"; -- Line 187   Column 6   Coefficient 0.00000000
         when "101110100110" => A <= "111111011001111001"; -- Line 187   Column 7   Coefficient -0.00930405
         when "101110100111" => A <= "000010011110111100"; -- Line 187   Column 8   Coefficient 0.03880310
         when "101110101000" => A <= "001111100101110011"; -- Line 187   Column 9   Coefficient 0.24360275
         when "101110101001" => A <= "111101111110110001"; -- Line 187   Column 10   Coefficient -0.03155136
         when "101110101010" => A <= "000000100001110011"; -- Line 187   Column 11   Coefficient 0.00825119
         when "101110101011" => A <= "000000000000110011"; -- Line 187   Column 12   Coefficient 0.00019455
         when "101110101100" => A <= "000000000000000000"; -- Line 187   Column 13   Coefficient 0.00000000
         when "101110101101" => A <= "000000000000000000"; -- Line 187   Column 14   Coefficient 0.00000000
         when "101110101110" => A <= "000000000000000000"; -- Line 187   Column 15   Coefficient 0.00000000
         when "101110101111" => A <= "000000000000000000"; -- Line 187   Column 16   Coefficient 0.00000000
         when "101110110000" => A <= "000000000000000000"; -- Line 188   Column 1   Coefficient 0.00000000
         when "101110110001" => A <= "000000000000000000"; -- Line 188   Column 2   Coefficient 0.00000000
         when "101110110010" => A <= "000000000000000000"; -- Line 188   Column 3   Coefficient 0.00000000
         when "101110110011" => A <= "000000000000000000"; -- Line 188   Column 4   Coefficient 0.00000000
         when "101110110100" => A <= "000000000000000000"; -- Line 188   Column 5   Coefficient 0.00000000
         when "101110110101" => A <= "000000000000000000"; -- Line 188   Column 6   Coefficient 0.00000000
         when "101110110110" => A <= "111111110001010101"; -- Line 188   Column 7   Coefficient -0.00358200
         when "101110110111" => A <= "000000100101011001"; -- Line 188   Column 8   Coefficient 0.00912857
         when "101110111000" => A <= "010001011110001011"; -- Line 188   Column 9   Coefficient 0.27299118
         when "101110111001" => A <= "111101011101101101"; -- Line 188   Column 10   Coefficient -0.03962326
         when "101110111010" => A <= "000000101011110101"; -- Line 188   Column 11   Coefficient 0.01070023
         when "101110111011" => A <= "000000000001100101"; -- Line 188   Column 12   Coefficient 0.00038528
         when "101110111100" => A <= "000000000000000000"; -- Line 188   Column 13   Coefficient 0.00000000
         when "101110111101" => A <= "000000000000000000"; -- Line 188   Column 14   Coefficient 0.00000000
         when "101110111110" => A <= "000000000000000000"; -- Line 188   Column 15   Coefficient 0.00000000
         when "101110111111" => A <= "000000000000000000"; -- Line 188   Column 16   Coefficient 0.00000000
         when "101111000000" => A <= "000000000000000000"; -- Line 189   Column 1   Coefficient 0.00000000
         when "101111000001" => A <= "000000000000000000"; -- Line 189   Column 2   Coefficient 0.00000000
         when "101111000010" => A <= "000000000000000000"; -- Line 189   Column 3   Coefficient 0.00000000
         when "101111000011" => A <= "000000000000000000"; -- Line 189   Column 4   Coefficient 0.00000000
         when "101111000100" => A <= "000000000000000000"; -- Line 189   Column 5   Coefficient 0.00000000
         when "101111000101" => A <= "000000000000000000"; -- Line 189   Column 6   Coefficient 0.00000000
         when "101111000110" => A <= "000000000111011010"; -- Line 189   Column 7   Coefficient 0.00180817
         when "101111000111" => A <= "111110110101100100"; -- Line 189   Column 8   Coefficient -0.01817322
         when "101111001000" => A <= "010011000101100111"; -- Line 189   Column 9   Coefficient 0.29824448
         when "101111001001" => A <= "111101000110110001"; -- Line 189   Column 10   Coefficient -0.04522324
         when "101111001010" => A <= "000000110100010110"; -- Line 189   Column 11   Coefficient 0.01277924
         when "101111001011" => A <= "000000000010010101"; -- Line 189   Column 12   Coefficient 0.00056839
         when "101111001100" => A <= "000000000000000000"; -- Line 189   Column 13   Coefficient 0.00000000
         when "101111001101" => A <= "000000000000000000"; -- Line 189   Column 14   Coefficient 0.00000000
         when "101111001110" => A <= "000000000000000000"; -- Line 189   Column 15   Coefficient 0.00000000
         when "101111001111" => A <= "000000000000000000"; -- Line 189   Column 16   Coefficient 0.00000000
         when "101111010000" => A <= "000000000000000000"; -- Line 190   Column 1   Coefficient 0.00000000
         when "101111010001" => A <= "000000000000000000"; -- Line 190   Column 2   Coefficient 0.00000000
         when "101111010010" => A <= "000000000000000000"; -- Line 190   Column 3   Coefficient 0.00000000
         when "101111010011" => A <= "000000000000000000"; -- Line 190   Column 4   Coefficient 0.00000000
         when "101111010100" => A <= "000000000000000000"; -- Line 190   Column 5   Coefficient 0.00000000
         when "101111010101" => A <= "000000000000000000"; -- Line 190   Column 6   Coefficient 0.00000000
         when "101111010110" => A <= "000000001111000010"; -- Line 190   Column 7   Coefficient 0.00366974
         when "101111010111" => A <= "111110000010011110"; -- Line 190   Column 8   Coefficient -0.03064728
         when "101111011000" => A <= "010011010010100110"; -- Line 190   Column 9   Coefficient 0.30141449
         when "101111011001" => A <= "111101100111001110"; -- Line 190   Column 10   Coefficient -0.03730011
         when "101111011010" => A <= "000000110010101110"; -- Line 190   Column 11   Coefficient 0.01238251
         when "101111011011" => A <= "000000000001111110"; -- Line 190   Column 12   Coefficient 0.00048065
         when "101111011100" => A <= "000000000000000000"; -- Line 190   Column 13   Coefficient 0.00000000
         when "101111011101" => A <= "000000000000000000"; -- Line 190   Column 14   Coefficient 0.00000000
         when "101111011110" => A <= "000000000000000000"; -- Line 190   Column 15   Coefficient 0.00000000
         when "101111011111" => A <= "000000000000000000"; -- Line 190   Column 16   Coefficient 0.00000000
         when "101111100000" => A <= "000000000000000000"; -- Line 191   Column 1   Coefficient 0.00000000
         when "101111100001" => A <= "000000000000000000"; -- Line 191   Column 2   Coefficient 0.00000000
         when "101111100010" => A <= "000000000000000000"; -- Line 191   Column 3   Coefficient 0.00000000
         when "101111100011" => A <= "000000000000000000"; -- Line 191   Column 4   Coefficient 0.00000000
         when "101111100100" => A <= "000000000000000000"; -- Line 191   Column 5   Coefficient 0.00000000
         when "101111100101" => A <= "000000000000000000"; -- Line 191   Column 6   Coefficient 0.00000000
         when "101111100110" => A <= "000000010000011000"; -- Line 191   Column 7   Coefficient 0.00399780
         when "101111100111" => A <= "111101101011101110"; -- Line 191   Column 8   Coefficient -0.03620148
         when "101111101000" => A <= "010010110100110100"; -- Line 191   Column 9   Coefficient 0.29414368
         when "101111101001" => A <= "111110100000101100"; -- Line 191   Column 10   Coefficient -0.02326965
         when "101111101010" => A <= "000000101101010111"; -- Line 191   Column 11   Coefficient 0.01107407
         when "101111101011" => A <= "000000000001000010"; -- Line 191   Column 12   Coefficient 0.00025177
         when "101111101100" => A <= "000000000000000000"; -- Line 191   Column 13   Coefficient 0.00000000
         when "101111101101" => A <= "000000000000000000"; -- Line 191   Column 14   Coefficient 0.00000000
         when "101111101110" => A <= "000000000000000000"; -- Line 191   Column 15   Coefficient 0.00000000
         when "101111101111" => A <= "000000000000000000"; -- Line 191   Column 16   Coefficient 0.00000000
         when "101111110000" => A <= "000000000000000000"; -- Line 192   Column 1   Coefficient 0.00000000
         when "101111110001" => A <= "000000000000000000"; -- Line 192   Column 2   Coefficient 0.00000000
         when "101111110010" => A <= "000000000000000000"; -- Line 192   Column 3   Coefficient 0.00000000
         when "101111110011" => A <= "000000000000000000"; -- Line 192   Column 4   Coefficient 0.00000000
         when "101111110100" => A <= "000000000000000000"; -- Line 192   Column 5   Coefficient 0.00000000
         when "101111110101" => A <= "000000000000000000"; -- Line 192   Column 6   Coefficient 0.00000000
         when "101111110110" => A <= "000000001111111100"; -- Line 192   Column 7   Coefficient 0.00389099
         when "101111110111" => A <= "111101100000101101"; -- Line 192   Column 8   Coefficient -0.03889084
         when "101111111000" => A <= "010010000001100011"; -- Line 192   Column 9   Coefficient 0.28162766
         when "101111111001" => A <= "111111101010001000"; -- Line 192   Column 10   Coefficient -0.00534058
         when "101111111010" => A <= "000000100010100100"; -- Line 192   Column 11   Coefficient 0.00843811
         when "101111111011" => A <= "000000000001001000"; -- Line 192   Column 12   Coefficient 0.00027466
         when "101111111100" => A <= "000000000000000000"; -- Line 192   Column 13   Coefficient 0.00000000
         when "101111111101" => A <= "000000000000000000"; -- Line 192   Column 14   Coefficient 0.00000000
         when "101111111110" => A <= "000000000000000000"; -- Line 192   Column 15   Coefficient 0.00000000
         when "101111111111" => A <= "000000000000000000"; -- Line 192   Column 16   Coefficient 0.00000000
         when "110000000000" => A <= "000000000000000000"; -- Line 193   Column 1   Coefficient 0.00000000
         when "110000000001" => A <= "000000000000000000"; -- Line 193   Column 2   Coefficient 0.00000000
         when "110000000010" => A <= "000000000000000000"; -- Line 193   Column 3   Coefficient 0.00000000
         when "110000000011" => A <= "000000000000000000"; -- Line 193   Column 4   Coefficient 0.00000000
         when "110000000100" => A <= "000000000000000000"; -- Line 193   Column 5   Coefficient 0.00000000
         when "110000000101" => A <= "000000000000000000"; -- Line 193   Column 6   Coefficient 0.00000000
         when "110000000110" => A <= "000000001101001100"; -- Line 193   Column 7   Coefficient 0.00321960
         when "110000000111" => A <= "111101100010001110"; -- Line 193   Column 8   Coefficient -0.03852081
         when "110000001000" => A <= "010000111010100101"; -- Line 193   Column 9   Coefficient 0.26430130
         when "110000001001" => A <= "000000111110100110"; -- Line 193   Column 10   Coefficient 0.01528168
         when "110000001010" => A <= "000000010110010000"; -- Line 193   Column 11   Coefficient 0.00543213
         when "110000001011" => A <= "000000000001001011"; -- Line 193   Column 12   Coefficient 0.00028610
         when "110000001100" => A <= "000000000000000000"; -- Line 193   Column 13   Coefficient 0.00000000
         when "110000001101" => A <= "000000000000000000"; -- Line 193   Column 14   Coefficient 0.00000000
         when "110000001110" => A <= "000000000000000000"; -- Line 193   Column 15   Coefficient 0.00000000
         when "110000001111" => A <= "000000000000000000"; -- Line 193   Column 16   Coefficient 0.00000000
         when "110000010000" => A <= "000000000000000000"; -- Line 194   Column 1   Coefficient 0.00000000
         when "110000010001" => A <= "000000000000000000"; -- Line 194   Column 2   Coefficient 0.00000000
         when "110000010010" => A <= "000000000000000000"; -- Line 194   Column 3   Coefficient 0.00000000
         when "110000010011" => A <= "000000000000000000"; -- Line 194   Column 4   Coefficient 0.00000000
         when "110000010100" => A <= "000000000000000000"; -- Line 194   Column 5   Coefficient 0.00000000
         when "110000010101" => A <= "000000000000000000"; -- Line 194   Column 6   Coefficient 0.00000000
         when "110000010110" => A <= "000000001010110110"; -- Line 194   Column 7   Coefficient 0.00264740
         when "110000010111" => A <= "111101100010101111"; -- Line 194   Column 8   Coefficient -0.03839493
         when "110000011000" => A <= "001111111010100001"; -- Line 194   Column 9   Coefficient 0.24866104
         when "110000011001" => A <= "000010000100001011"; -- Line 194   Column 10   Coefficient 0.03226852
         when "110000011010" => A <= "000000010100110111"; -- Line 194   Column 11   Coefficient 0.00509262
         when "110000011011" => A <= "111111111110110111"; -- Line 194   Column 12   Coefficient -0.00027847
         when "110000011100" => A <= "000000000000000000"; -- Line 194   Column 13   Coefficient 0.00000000
         when "110000011101" => A <= "000000000000000000"; -- Line 194   Column 14   Coefficient 0.00000000
         when "110000011110" => A <= "000000000000000000"; -- Line 194   Column 15   Coefficient 0.00000000
         when "110000011111" => A <= "000000000000000000"; -- Line 194   Column 16   Coefficient 0.00000000
         when "110000100000" => A <= "000000000000000000"; -- Line 195   Column 1   Coefficient 0.00000000
         when "110000100001" => A <= "000000000000000000"; -- Line 195   Column 2   Coefficient 0.00000000
         when "110000100010" => A <= "000000000000000000"; -- Line 195   Column 3   Coefficient 0.00000000
         when "110000100011" => A <= "000000000000000000"; -- Line 195   Column 4   Coefficient 0.00000000
         when "110000100100" => A <= "000000000000000000"; -- Line 195   Column 5   Coefficient 0.00000000
         when "110000100101" => A <= "000000000000000000"; -- Line 195   Column 6   Coefficient 0.00000000
         when "110000100110" => A <= "000000001000010011"; -- Line 195   Column 7   Coefficient 0.00202560
         when "110000100111" => A <= "111101100110110000"; -- Line 195   Column 8   Coefficient -0.03741455
         when "110000101000" => A <= "001110110101010100"; -- Line 195   Column 9   Coefficient 0.23176575
         when "110000101001" => A <= "000011001010010011"; -- Line 195   Column 10   Coefficient 0.04938889
         when "110000101010" => A <= "000000010100111001"; -- Line 195   Column 11   Coefficient 0.00510025
         when "110000101011" => A <= "111111111100011110"; -- Line 195   Column 12   Coefficient -0.00086212
         when "110000101100" => A <= "111111111111111111"; -- Line 195   Column 13   Coefficient -0.00000381
         when "110000101101" => A <= "000000000000000000"; -- Line 195   Column 14   Coefficient 0.00000000
         when "110000101110" => A <= "000000000000000000"; -- Line 195   Column 15   Coefficient 0.00000000
         when "110000101111" => A <= "000000000000000000"; -- Line 195   Column 16   Coefficient 0.00000000
         when "110000110000" => A <= "000000000000000000"; -- Line 196   Column 1   Coefficient 0.00000000
         when "110000110001" => A <= "000000000000000000"; -- Line 196   Column 2   Coefficient 0.00000000
         when "110000110010" => A <= "000000000000000000"; -- Line 196   Column 3   Coefficient 0.00000000
         when "110000110011" => A <= "000000000000000000"; -- Line 196   Column 4   Coefficient 0.00000000
         when "110000110100" => A <= "000000000000000000"; -- Line 196   Column 5   Coefficient 0.00000000
         when "110000110101" => A <= "000000000000000000"; -- Line 196   Column 6   Coefficient 0.00000000
         when "110000110110" => A <= "000000000011111000"; -- Line 196   Column 7   Coefficient 0.00094604
         when "110000110111" => A <= "111101110100001010"; -- Line 196   Column 8   Coefficient -0.03414154
         when "110000111000" => A <= "001101100011111111"; -- Line 196   Column 9   Coefficient 0.21191025
         when "110000111001" => A <= "000100010011001101"; -- Line 196   Column 10   Coefficient 0.06718826
         when "110000111010" => A <= "000000010111101010"; -- Line 196   Column 11   Coefficient 0.00577545
         when "110000111011" => A <= "111111111001000110"; -- Line 196   Column 12   Coefficient -0.00168610
         when "110000111100" => A <= "000000000000000011"; -- Line 196   Column 13   Coefficient 0.00001144
         when "110000111101" => A <= "000000000000000000"; -- Line 196   Column 14   Coefficient 0.00000000
         when "110000111110" => A <= "000000000000000000"; -- Line 196   Column 15   Coefficient 0.00000000
         when "110000111111" => A <= "000000000000000000"; -- Line 196   Column 16   Coefficient 0.00000000
         when "110001000000" => A <= "000000000000000000"; -- Line 197   Column 1   Coefficient 0.00000000
         when "110001000001" => A <= "000000000000000000"; -- Line 197   Column 2   Coefficient 0.00000000
         when "110001000010" => A <= "000000000000000000"; -- Line 197   Column 3   Coefficient 0.00000000
         when "110001000011" => A <= "000000000000000000"; -- Line 197   Column 4   Coefficient 0.00000000
         when "110001000100" => A <= "000000000000000000"; -- Line 197   Column 5   Coefficient 0.00000000
         when "110001000101" => A <= "000000000000000000"; -- Line 197   Column 6   Coefficient 0.00000000
         when "110001000110" => A <= "111111111111010011"; -- Line 197   Column 7   Coefficient -0.00017166
         when "110001000111" => A <= "111110000101010011"; -- Line 197   Column 8   Coefficient -0.02995682
         when "110001001000" => A <= "001100001011101000"; -- Line 197   Column 9   Coefficient 0.19033813
         when "110001001001" => A <= "000101100000010101"; -- Line 197   Column 10   Coefficient 0.08601761
         when "110001001010" => A <= "000000011000110111"; -- Line 197   Column 11   Coefficient 0.00606918
         when "110001001011" => A <= "111111110110011111"; -- Line 197   Column 12   Coefficient -0.00232315
         when "110001001100" => A <= "000000000000000110"; -- Line 197   Column 13   Coefficient 0.00002289
         when "110001001101" => A <= "000000000000000000"; -- Line 197   Column 14   Coefficient 0.00000000
         when "110001001110" => A <= "000000000000000000"; -- Line 197   Column 15   Coefficient 0.00000000
         when "110001001111" => A <= "000000000000000000"; -- Line 197   Column 16   Coefficient 0.00000000
         when "110001010000" => A <= "000000000000000000"; -- Line 198   Column 1   Coefficient 0.00000000
         when "110001010001" => A <= "000000000000000000"; -- Line 198   Column 2   Coefficient 0.00000000
         when "110001010010" => A <= "000000000000000000"; -- Line 198   Column 3   Coefficient 0.00000000
         when "110001010011" => A <= "000000000000000000"; -- Line 198   Column 4   Coefficient 0.00000000
         when "110001010100" => A <= "000000000000000000"; -- Line 198   Column 5   Coefficient 0.00000000
         when "110001010101" => A <= "000000000000000000"; -- Line 198   Column 6   Coefficient 0.00000000
         when "110001010110" => A <= "111111111110010010"; -- Line 198   Column 7   Coefficient -0.00041962
         when "110001010111" => A <= "111110010000110000"; -- Line 198   Column 8   Coefficient -0.02716064
         when "110001011000" => A <= "001010101100000111"; -- Line 198   Column 9   Coefficient 0.16701889
         when "110001011001" => A <= "000111000101010101"; -- Line 198   Column 10   Coefficient 0.11067581
         when "110001011010" => A <= "000000000100100100"; -- Line 198   Column 11   Coefficient 0.00111389
         when "110001011011" => A <= "111111111010111001"; -- Line 198   Column 12   Coefficient -0.00124741
         when "110001011100" => A <= "000000000000000100"; -- Line 198   Column 13   Coefficient 0.00001526
         when "110001011101" => A <= "000000000000000000"; -- Line 198   Column 14   Coefficient 0.00000000
         when "110001011110" => A <= "000000000000000000"; -- Line 198   Column 15   Coefficient 0.00000000
         when "110001011111" => A <= "000000000000000000"; -- Line 198   Column 16   Coefficient 0.00000000
         when "110001100000" => A <= "000000000000000000"; -- Line 199   Column 1   Coefficient 0.00000000
         when "110001100001" => A <= "000000000000000000"; -- Line 199   Column 2   Coefficient 0.00000000
         when "110001100010" => A <= "000000000000000000"; -- Line 199   Column 3   Coefficient 0.00000000
         when "110001100011" => A <= "000000000000000000"; -- Line 199   Column 4   Coefficient 0.00000000
         when "110001100100" => A <= "000000000000000000"; -- Line 199   Column 5   Coefficient 0.00000000
         when "110001100101" => A <= "000000000000000000"; -- Line 199   Column 6   Coefficient 0.00000000
         when "110001100110" => A <= "111111111110100110"; -- Line 199   Column 7   Coefficient -0.00034332
         when "110001100111" => A <= "111110011011111010"; -- Line 199   Column 8   Coefficient -0.02443695
         when "110001101000" => A <= "001001000110101001"; -- Line 199   Column 9   Coefficient 0.14224625
         when "110001101001" => A <= "001000110101000000"; -- Line 199   Column 10   Coefficient 0.13793945
         when "110001101010" => A <= "111111100111100010"; -- Line 199   Column 11   Coefficient -0.00597382
         when "110001101011" => A <= "000000000010010011"; -- Line 199   Column 12   Coefficient 0.00056076
         when "110001101100" => A <= "000000000000000011"; -- Line 199   Column 13   Coefficient 0.00001144
         when "110001101101" => A <= "000000000000000000"; -- Line 199   Column 14   Coefficient 0.00000000
         when "110001101110" => A <= "000000000000000000"; -- Line 199   Column 15   Coefficient 0.00000000
         when "110001101111" => A <= "000000000000000000"; -- Line 199   Column 16   Coefficient 0.00000000
         when "110001110000" => A <= "000000000000000000"; -- Line 200   Column 1   Coefficient 0.00000000
         when "110001110001" => A <= "000000000000000000"; -- Line 200   Column 2   Coefficient 0.00000000
         when "110001110010" => A <= "000000000000000000"; -- Line 200   Column 3   Coefficient 0.00000000
         when "110001110011" => A <= "000000000000000000"; -- Line 200   Column 4   Coefficient 0.00000000
         when "110001110100" => A <= "000000000000000000"; -- Line 200   Column 5   Coefficient 0.00000000
         when "110001110101" => A <= "000000000000000000"; -- Line 200   Column 6   Coefficient 0.00000000
         when "110001110110" => A <= "111111111111001011"; -- Line 200   Column 7   Coefficient -0.00020218
         when "110001110111" => A <= "111110100110010011"; -- Line 200   Column 8   Coefficient -0.02190018
         when "110001111000" => A <= "000111100110110001"; -- Line 200   Column 9   Coefficient 0.11883926
         when "110001111001" => A <= "001010011001111000"; -- Line 200   Column 10   Coefficient 0.16256714
         when "110001111010" => A <= "111111010000101110"; -- Line 200   Column 11   Coefficient -0.01154327
         when "110001111011" => A <= "000000001001011000"; -- Line 200   Column 12   Coefficient 0.00228882
         when "110001111100" => A <= "111111111111110100"; -- Line 200   Column 13   Coefficient -0.00004578
         when "110001111101" => A <= "000000000000000000"; -- Line 200   Column 14   Coefficient 0.00000000
         when "110001111110" => A <= "000000000000000000"; -- Line 200   Column 15   Coefficient 0.00000000
         when "110001111111" => A <= "000000000000000000"; -- Line 200   Column 16   Coefficient 0.00000000
         when "110010000000" => A <= "000000000000000000"; -- Line 201   Column 1   Coefficient 0.00000000
         when "110010000001" => A <= "000000000000000000"; -- Line 201   Column 2   Coefficient 0.00000000
         when "110010000010" => A <= "000000000000000000"; -- Line 201   Column 3   Coefficient 0.00000000
         when "110010000011" => A <= "000000000000000000"; -- Line 201   Column 4   Coefficient 0.00000000
         when "110010000100" => A <= "000000000000000000"; -- Line 201   Column 5   Coefficient 0.00000000
         when "110010000101" => A <= "000000000000000000"; -- Line 201   Column 6   Coefficient 0.00000000
         when "110010000110" => A <= "000000000000000011"; -- Line 201   Column 7   Coefficient 0.00001144
         when "110010000111" => A <= "111110110001100001"; -- Line 201   Column 8   Coefficient -0.01916122
         when "110010001000" => A <= "000110000101110011"; -- Line 201   Column 9   Coefficient 0.09516525
         when "110010001001" => A <= "001011111101111010"; -- Line 201   Column 10   Coefficient 0.18698883
         when "110010001010" => A <= "111110111010000001"; -- Line 201   Column 11   Coefficient -0.01708603
         when "110010001011" => A <= "000000010001001000"; -- Line 201   Column 12   Coefficient 0.00418091
         when "110010001100" => A <= "111111111111100110"; -- Line 201   Column 13   Coefficient -0.00009918
         when "110010001101" => A <= "000000000000000000"; -- Line 201   Column 14   Coefficient 0.00000000
         when "110010001110" => A <= "000000000000000000"; -- Line 201   Column 15   Coefficient 0.00000000
         when "110010001111" => A <= "000000000000000000"; -- Line 201   Column 16   Coefficient 0.00000000
         when "110010010000" => A <= "000000000000000000"; -- Line 202   Column 1   Coefficient 0.00000000
         when "110010010001" => A <= "000000000000000000"; -- Line 202   Column 2   Coefficient 0.00000000
         when "110010010010" => A <= "000000000000000000"; -- Line 202   Column 3   Coefficient 0.00000000
         when "110010010011" => A <= "000000000000000000"; -- Line 202   Column 4   Coefficient 0.00000000
         when "110010010100" => A <= "000000000000000000"; -- Line 202   Column 5   Coefficient 0.00000000
         when "110010010101" => A <= "000000000000000000"; -- Line 202   Column 6   Coefficient 0.00000000
         when "110010010110" => A <= "000000000000001001"; -- Line 202   Column 7   Coefficient 0.00003433
         when "110010010111" => A <= "111111000100111001"; -- Line 202   Column 8   Coefficient -0.01443100
         when "110010011000" => A <= "000100010010000101"; -- Line 202   Column 9   Coefficient 0.06691360
         when "110010011001" => A <= "001101110100101001"; -- Line 202   Column 10   Coefficient 0.21597672
         when "110010011010" => A <= "111110011010010101"; -- Line 202   Column 11   Coefficient -0.02482224
         when "110010011011" => A <= "000000011001110100"; -- Line 202   Column 12   Coefficient 0.00630188
         when "110010011100" => A <= "000000000000000111"; -- Line 202   Column 13   Coefficient 0.00002670
         when "110010011101" => A <= "000000000000000000"; -- Line 202   Column 14   Coefficient 0.00000000
         when "110010011110" => A <= "000000000000000000"; -- Line 202   Column 15   Coefficient 0.00000000
         when "110010011111" => A <= "000000000000000000"; -- Line 202   Column 16   Coefficient 0.00000000
         when "110010100000" => A <= "000000000000000000"; -- Line 203   Column 1   Coefficient 0.00000000
         when "110010100001" => A <= "000000000000000000"; -- Line 203   Column 2   Coefficient 0.00000000
         when "110010100010" => A <= "000000000000000000"; -- Line 203   Column 3   Coefficient 0.00000000
         when "110010100011" => A <= "000000000000000000"; -- Line 203   Column 4   Coefficient 0.00000000
         when "110010100100" => A <= "000000000000000000"; -- Line 203   Column 5   Coefficient 0.00000000
         when "110010100101" => A <= "000000000000000000"; -- Line 203   Column 6   Coefficient 0.00000000
         when "110010100110" => A <= "000000000000000000"; -- Line 203   Column 7   Coefficient 0.00000000
         when "110010100111" => A <= "111111011001111001"; -- Line 203   Column 8   Coefficient -0.00930405
         when "110010101000" => A <= "000010011110111100"; -- Line 203   Column 9   Coefficient 0.03880310
         when "110010101001" => A <= "001111100101110011"; -- Line 203   Column 10   Coefficient 0.24360275
         when "110010101010" => A <= "111101111110110001"; -- Line 203   Column 11   Coefficient -0.03155136
         when "110010101011" => A <= "000000100001110011"; -- Line 203   Column 12   Coefficient 0.00825119
         when "110010101100" => A <= "000000000000110011"; -- Line 203   Column 13   Coefficient 0.00019455
         when "110010101101" => A <= "000000000000000000"; -- Line 203   Column 14   Coefficient 0.00000000
         when "110010101110" => A <= "000000000000000000"; -- Line 203   Column 15   Coefficient 0.00000000
         when "110010101111" => A <= "000000000000000000"; -- Line 203   Column 16   Coefficient 0.00000000
         when "110010110000" => A <= "000000000000000000"; -- Line 204   Column 1   Coefficient 0.00000000
         when "110010110001" => A <= "000000000000000000"; -- Line 204   Column 2   Coefficient 0.00000000
         when "110010110010" => A <= "000000000000000000"; -- Line 204   Column 3   Coefficient 0.00000000
         when "110010110011" => A <= "000000000000000000"; -- Line 204   Column 4   Coefficient 0.00000000
         when "110010110100" => A <= "000000000000000000"; -- Line 204   Column 5   Coefficient 0.00000000
         when "110010110101" => A <= "000000000000000000"; -- Line 204   Column 6   Coefficient 0.00000000
         when "110010110110" => A <= "000000000000000000"; -- Line 204   Column 7   Coefficient 0.00000000
         when "110010110111" => A <= "111111110001010101"; -- Line 204   Column 8   Coefficient -0.00358200
         when "110010111000" => A <= "000000100101011001"; -- Line 204   Column 9   Coefficient 0.00912857
         when "110010111001" => A <= "010001011110001011"; -- Line 204   Column 10   Coefficient 0.27299118
         when "110010111010" => A <= "111101011101101101"; -- Line 204   Column 11   Coefficient -0.03962326
         when "110010111011" => A <= "000000101011110101"; -- Line 204   Column 12   Coefficient 0.01070023
         when "110010111100" => A <= "000000000001100101"; -- Line 204   Column 13   Coefficient 0.00038528
         when "110010111101" => A <= "000000000000000000"; -- Line 204   Column 14   Coefficient 0.00000000
         when "110010111110" => A <= "000000000000000000"; -- Line 204   Column 15   Coefficient 0.00000000
         when "110010111111" => A <= "000000000000000000"; -- Line 204   Column 16   Coefficient 0.00000000
         when "110011000000" => A <= "000000000000000000"; -- Line 205   Column 1   Coefficient 0.00000000
         when "110011000001" => A <= "000000000000000000"; -- Line 205   Column 2   Coefficient 0.00000000
         when "110011000010" => A <= "000000000000000000"; -- Line 205   Column 3   Coefficient 0.00000000
         when "110011000011" => A <= "000000000000000000"; -- Line 205   Column 4   Coefficient 0.00000000
         when "110011000100" => A <= "000000000000000000"; -- Line 205   Column 5   Coefficient 0.00000000
         when "110011000101" => A <= "000000000000000000"; -- Line 205   Column 6   Coefficient 0.00000000
         when "110011000110" => A <= "000000000000000000"; -- Line 205   Column 7   Coefficient 0.00000000
         when "110011000111" => A <= "000000000111011010"; -- Line 205   Column 8   Coefficient 0.00180817
         when "110011001000" => A <= "111110110101100100"; -- Line 205   Column 9   Coefficient -0.01817322
         when "110011001001" => A <= "010011000101100111"; -- Line 205   Column 10   Coefficient 0.29824448
         when "110011001010" => A <= "111101000110110001"; -- Line 205   Column 11   Coefficient -0.04522324
         when "110011001011" => A <= "000000110100010110"; -- Line 205   Column 12   Coefficient 0.01277924
         when "110011001100" => A <= "000000000010010101"; -- Line 205   Column 13   Coefficient 0.00056839
         when "110011001101" => A <= "000000000000000000"; -- Line 205   Column 14   Coefficient 0.00000000
         when "110011001110" => A <= "000000000000000000"; -- Line 205   Column 15   Coefficient 0.00000000
         when "110011001111" => A <= "000000000000000000"; -- Line 205   Column 16   Coefficient 0.00000000
         when "110011010000" => A <= "000000000000000000"; -- Line 206   Column 1   Coefficient 0.00000000
         when "110011010001" => A <= "000000000000000000"; -- Line 206   Column 2   Coefficient 0.00000000
         when "110011010010" => A <= "000000000000000000"; -- Line 206   Column 3   Coefficient 0.00000000
         when "110011010011" => A <= "000000000000000000"; -- Line 206   Column 4   Coefficient 0.00000000
         when "110011010100" => A <= "000000000000000000"; -- Line 206   Column 5   Coefficient 0.00000000
         when "110011010101" => A <= "000000000000000000"; -- Line 206   Column 6   Coefficient 0.00000000
         when "110011010110" => A <= "000000000000000000"; -- Line 206   Column 7   Coefficient 0.00000000
         when "110011010111" => A <= "000000001111000010"; -- Line 206   Column 8   Coefficient 0.00366974
         when "110011011000" => A <= "111110000010011110"; -- Line 206   Column 9   Coefficient -0.03064728
         when "110011011001" => A <= "010011010010100110"; -- Line 206   Column 10   Coefficient 0.30141449
         when "110011011010" => A <= "111101100111001110"; -- Line 206   Column 11   Coefficient -0.03730011
         when "110011011011" => A <= "000000110010101110"; -- Line 206   Column 12   Coefficient 0.01238251
         when "110011011100" => A <= "000000000001111110"; -- Line 206   Column 13   Coefficient 0.00048065
         when "110011011101" => A <= "000000000000000000"; -- Line 206   Column 14   Coefficient 0.00000000
         when "110011011110" => A <= "000000000000000000"; -- Line 206   Column 15   Coefficient 0.00000000
         when "110011011111" => A <= "000000000000000000"; -- Line 206   Column 16   Coefficient 0.00000000
         when "110011100000" => A <= "000000000000000000"; -- Line 207   Column 1   Coefficient 0.00000000
         when "110011100001" => A <= "000000000000000000"; -- Line 207   Column 2   Coefficient 0.00000000
         when "110011100010" => A <= "000000000000000000"; -- Line 207   Column 3   Coefficient 0.00000000
         when "110011100011" => A <= "000000000000000000"; -- Line 207   Column 4   Coefficient 0.00000000
         when "110011100100" => A <= "000000000000000000"; -- Line 207   Column 5   Coefficient 0.00000000
         when "110011100101" => A <= "000000000000000000"; -- Line 207   Column 6   Coefficient 0.00000000
         when "110011100110" => A <= "000000000000000000"; -- Line 207   Column 7   Coefficient 0.00000000
         when "110011100111" => A <= "000000010000011000"; -- Line 207   Column 8   Coefficient 0.00399780
         when "110011101000" => A <= "111101101011101110"; -- Line 207   Column 9   Coefficient -0.03620148
         when "110011101001" => A <= "010010110100110100"; -- Line 207   Column 10   Coefficient 0.29414368
         when "110011101010" => A <= "111110100000101100"; -- Line 207   Column 11   Coefficient -0.02326965
         when "110011101011" => A <= "000000101101010111"; -- Line 207   Column 12   Coefficient 0.01107407
         when "110011101100" => A <= "000000000001000010"; -- Line 207   Column 13   Coefficient 0.00025177
         when "110011101101" => A <= "000000000000000000"; -- Line 207   Column 14   Coefficient 0.00000000
         when "110011101110" => A <= "000000000000000000"; -- Line 207   Column 15   Coefficient 0.00000000
         when "110011101111" => A <= "000000000000000000"; -- Line 207   Column 16   Coefficient 0.00000000
         when "110011110000" => A <= "000000000000000000"; -- Line 208   Column 1   Coefficient 0.00000000
         when "110011110001" => A <= "000000000000000000"; -- Line 208   Column 2   Coefficient 0.00000000
         when "110011110010" => A <= "000000000000000000"; -- Line 208   Column 3   Coefficient 0.00000000
         when "110011110011" => A <= "000000000000000000"; -- Line 208   Column 4   Coefficient 0.00000000
         when "110011110100" => A <= "000000000000000000"; -- Line 208   Column 5   Coefficient 0.00000000
         when "110011110101" => A <= "000000000000000000"; -- Line 208   Column 6   Coefficient 0.00000000
         when "110011110110" => A <= "000000000000000000"; -- Line 208   Column 7   Coefficient 0.00000000
         when "110011110111" => A <= "000000001111111100"; -- Line 208   Column 8   Coefficient 0.00389099
         when "110011111000" => A <= "111101100000101101"; -- Line 208   Column 9   Coefficient -0.03889084
         when "110011111001" => A <= "010010000001100011"; -- Line 208   Column 10   Coefficient 0.28162766
         when "110011111010" => A <= "111111101010001000"; -- Line 208   Column 11   Coefficient -0.00534058
         when "110011111011" => A <= "000000100010100100"; -- Line 208   Column 12   Coefficient 0.00843811
         when "110011111100" => A <= "000000000001001000"; -- Line 208   Column 13   Coefficient 0.00027466
         when "110011111101" => A <= "000000000000000000"; -- Line 208   Column 14   Coefficient 0.00000000
         when "110011111110" => A <= "000000000000000000"; -- Line 208   Column 15   Coefficient 0.00000000
         when "110011111111" => A <= "000000000000000000"; -- Line 208   Column 16   Coefficient 0.00000000
         when "110100000000" => A <= "000000000000000000"; -- Line 209   Column 1   Coefficient 0.00000000
         when "110100000001" => A <= "000000000000000000"; -- Line 209   Column 2   Coefficient 0.00000000
         when "110100000010" => A <= "000000000000000000"; -- Line 209   Column 3   Coefficient 0.00000000
         when "110100000011" => A <= "000000000000000000"; -- Line 209   Column 4   Coefficient 0.00000000
         when "110100000100" => A <= "000000000000000000"; -- Line 209   Column 5   Coefficient 0.00000000
         when "110100000101" => A <= "000000000000000000"; -- Line 209   Column 6   Coefficient 0.00000000
         when "110100000110" => A <= "000000000000000000"; -- Line 209   Column 7   Coefficient 0.00000000
         when "110100000111" => A <= "000000001101001100"; -- Line 209   Column 8   Coefficient 0.00321960
         when "110100001000" => A <= "111101100010001110"; -- Line 209   Column 9   Coefficient -0.03852081
         when "110100001001" => A <= "010000111010100101"; -- Line 209   Column 10   Coefficient 0.26430130
         when "110100001010" => A <= "000000111110100110"; -- Line 209   Column 11   Coefficient 0.01528168
         when "110100001011" => A <= "000000010110010000"; -- Line 209   Column 12   Coefficient 0.00543213
         when "110100001100" => A <= "000000000001001011"; -- Line 209   Column 13   Coefficient 0.00028610
         when "110100001101" => A <= "000000000000000000"; -- Line 209   Column 14   Coefficient 0.00000000
         when "110100001110" => A <= "000000000000000000"; -- Line 209   Column 15   Coefficient 0.00000000
         when "110100001111" => A <= "000000000000000000"; -- Line 209   Column 16   Coefficient 0.00000000
         when "110100010000" => A <= "000000000000000000"; -- Line 210   Column 1   Coefficient 0.00000000
         when "110100010001" => A <= "000000000000000000"; -- Line 210   Column 2   Coefficient 0.00000000
         when "110100010010" => A <= "000000000000000000"; -- Line 210   Column 3   Coefficient 0.00000000
         when "110100010011" => A <= "000000000000000000"; -- Line 210   Column 4   Coefficient 0.00000000
         when "110100010100" => A <= "000000000000000000"; -- Line 210   Column 5   Coefficient 0.00000000
         when "110100010101" => A <= "000000000000000000"; -- Line 210   Column 6   Coefficient 0.00000000
         when "110100010110" => A <= "000000000000000000"; -- Line 210   Column 7   Coefficient 0.00000000
         when "110100010111" => A <= "000000001010110110"; -- Line 210   Column 8   Coefficient 0.00264740
         when "110100011000" => A <= "111101100010101111"; -- Line 210   Column 9   Coefficient -0.03839493
         when "110100011001" => A <= "001111111010100001"; -- Line 210   Column 10   Coefficient 0.24866104
         when "110100011010" => A <= "000010000100001011"; -- Line 210   Column 11   Coefficient 0.03226852
         when "110100011011" => A <= "000000010100110111"; -- Line 210   Column 12   Coefficient 0.00509262
         when "110100011100" => A <= "111111111110110111"; -- Line 210   Column 13   Coefficient -0.00027847
         when "110100011101" => A <= "000000000000000000"; -- Line 210   Column 14   Coefficient 0.00000000
         when "110100011110" => A <= "000000000000000000"; -- Line 210   Column 15   Coefficient 0.00000000
         when "110100011111" => A <= "000000000000000000"; -- Line 210   Column 16   Coefficient 0.00000000
         when "110100100000" => A <= "000000000000000000"; -- Line 211   Column 1   Coefficient 0.00000000
         when "110100100001" => A <= "000000000000000000"; -- Line 211   Column 2   Coefficient 0.00000000
         when "110100100010" => A <= "000000000000000000"; -- Line 211   Column 3   Coefficient 0.00000000
         when "110100100011" => A <= "000000000000000000"; -- Line 211   Column 4   Coefficient 0.00000000
         when "110100100100" => A <= "000000000000000000"; -- Line 211   Column 5   Coefficient 0.00000000
         when "110100100101" => A <= "000000000000000000"; -- Line 211   Column 6   Coefficient 0.00000000
         when "110100100110" => A <= "000000000000000000"; -- Line 211   Column 7   Coefficient 0.00000000
         when "110100100111" => A <= "000000001000010011"; -- Line 211   Column 8   Coefficient 0.00202560
         when "110100101000" => A <= "111101100110110000"; -- Line 211   Column 9   Coefficient -0.03741455
         when "110100101001" => A <= "001110110101010100"; -- Line 211   Column 10   Coefficient 0.23176575
         when "110100101010" => A <= "000011001010010011"; -- Line 211   Column 11   Coefficient 0.04938889
         when "110100101011" => A <= "000000010100111001"; -- Line 211   Column 12   Coefficient 0.00510025
         when "110100101100" => A <= "111111111100011110"; -- Line 211   Column 13   Coefficient -0.00086212
         when "110100101101" => A <= "111111111111111111"; -- Line 211   Column 14   Coefficient -0.00000381
         when "110100101110" => A <= "000000000000000000"; -- Line 211   Column 15   Coefficient 0.00000000
         when "110100101111" => A <= "000000000000000000"; -- Line 211   Column 16   Coefficient 0.00000000
         when "110100110000" => A <= "000000000000000000"; -- Line 212   Column 1   Coefficient 0.00000000
         when "110100110001" => A <= "000000000000000000"; -- Line 212   Column 2   Coefficient 0.00000000
         when "110100110010" => A <= "000000000000000000"; -- Line 212   Column 3   Coefficient 0.00000000
         when "110100110011" => A <= "000000000000000000"; -- Line 212   Column 4   Coefficient 0.00000000
         when "110100110100" => A <= "000000000000000000"; -- Line 212   Column 5   Coefficient 0.00000000
         when "110100110101" => A <= "000000000000000000"; -- Line 212   Column 6   Coefficient 0.00000000
         when "110100110110" => A <= "000000000000000000"; -- Line 212   Column 7   Coefficient 0.00000000
         when "110100110111" => A <= "000000000011111000"; -- Line 212   Column 8   Coefficient 0.00094604
         when "110100111000" => A <= "111101110100001010"; -- Line 212   Column 9   Coefficient -0.03414154
         when "110100111001" => A <= "001101100011111111"; -- Line 212   Column 10   Coefficient 0.21191025
         when "110100111010" => A <= "000100010011001101"; -- Line 212   Column 11   Coefficient 0.06718826
         when "110100111011" => A <= "000000010111101010"; -- Line 212   Column 12   Coefficient 0.00577545
         when "110100111100" => A <= "111111111001000110"; -- Line 212   Column 13   Coefficient -0.00168610
         when "110100111101" => A <= "000000000000000011"; -- Line 212   Column 14   Coefficient 0.00001144
         when "110100111110" => A <= "000000000000000000"; -- Line 212   Column 15   Coefficient 0.00000000
         when "110100111111" => A <= "000000000000000000"; -- Line 212   Column 16   Coefficient 0.00000000
         when "110101000000" => A <= "000000000000000000"; -- Line 213   Column 1   Coefficient 0.00000000
         when "110101000001" => A <= "000000000000000000"; -- Line 213   Column 2   Coefficient 0.00000000
         when "110101000010" => A <= "000000000000000000"; -- Line 213   Column 3   Coefficient 0.00000000
         when "110101000011" => A <= "000000000000000000"; -- Line 213   Column 4   Coefficient 0.00000000
         when "110101000100" => A <= "000000000000000000"; -- Line 213   Column 5   Coefficient 0.00000000
         when "110101000101" => A <= "000000000000000000"; -- Line 213   Column 6   Coefficient 0.00000000
         when "110101000110" => A <= "000000000000000000"; -- Line 213   Column 7   Coefficient 0.00000000
         when "110101000111" => A <= "111111111111010011"; -- Line 213   Column 8   Coefficient -0.00017166
         when "110101001000" => A <= "111110000101010011"; -- Line 213   Column 9   Coefficient -0.02995682
         when "110101001001" => A <= "001100001011101000"; -- Line 213   Column 10   Coefficient 0.19033813
         when "110101001010" => A <= "000101100000010101"; -- Line 213   Column 11   Coefficient 0.08601761
         when "110101001011" => A <= "000000011000110111"; -- Line 213   Column 12   Coefficient 0.00606918
         when "110101001100" => A <= "111111110110011111"; -- Line 213   Column 13   Coefficient -0.00232315
         when "110101001101" => A <= "000000000000000110"; -- Line 213   Column 14   Coefficient 0.00002289
         when "110101001110" => A <= "000000000000000000"; -- Line 213   Column 15   Coefficient 0.00000000
         when "110101001111" => A <= "000000000000000000"; -- Line 213   Column 16   Coefficient 0.00000000
         when "110101010000" => A <= "000000000000000000"; -- Line 214   Column 1   Coefficient 0.00000000
         when "110101010001" => A <= "000000000000000000"; -- Line 214   Column 2   Coefficient 0.00000000
         when "110101010010" => A <= "000000000000000000"; -- Line 214   Column 3   Coefficient 0.00000000
         when "110101010011" => A <= "000000000000000000"; -- Line 214   Column 4   Coefficient 0.00000000
         when "110101010100" => A <= "000000000000000000"; -- Line 214   Column 5   Coefficient 0.00000000
         when "110101010101" => A <= "000000000000000000"; -- Line 214   Column 6   Coefficient 0.00000000
         when "110101010110" => A <= "000000000000000000"; -- Line 214   Column 7   Coefficient 0.00000000
         when "110101010111" => A <= "111111111110010010"; -- Line 214   Column 8   Coefficient -0.00041962
         when "110101011000" => A <= "111110010000110000"; -- Line 214   Column 9   Coefficient -0.02716064
         when "110101011001" => A <= "001010101100000111"; -- Line 214   Column 10   Coefficient 0.16701889
         when "110101011010" => A <= "000111000101010101"; -- Line 214   Column 11   Coefficient 0.11067581
         when "110101011011" => A <= "000000000100100100"; -- Line 214   Column 12   Coefficient 0.00111389
         when "110101011100" => A <= "111111111010111001"; -- Line 214   Column 13   Coefficient -0.00124741
         when "110101011101" => A <= "000000000000000100"; -- Line 214   Column 14   Coefficient 0.00001526
         when "110101011110" => A <= "000000000000000000"; -- Line 214   Column 15   Coefficient 0.00000000
         when "110101011111" => A <= "000000000000000000"; -- Line 214   Column 16   Coefficient 0.00000000
         when "110101100000" => A <= "000000000000000000"; -- Line 215   Column 1   Coefficient 0.00000000
         when "110101100001" => A <= "000000000000000000"; -- Line 215   Column 2   Coefficient 0.00000000
         when "110101100010" => A <= "000000000000000000"; -- Line 215   Column 3   Coefficient 0.00000000
         when "110101100011" => A <= "000000000000000000"; -- Line 215   Column 4   Coefficient 0.00000000
         when "110101100100" => A <= "000000000000000000"; -- Line 215   Column 5   Coefficient 0.00000000
         when "110101100101" => A <= "000000000000000000"; -- Line 215   Column 6   Coefficient 0.00000000
         when "110101100110" => A <= "000000000000000000"; -- Line 215   Column 7   Coefficient 0.00000000
         when "110101100111" => A <= "111111111110100110"; -- Line 215   Column 8   Coefficient -0.00034332
         when "110101101000" => A <= "111110011011111010"; -- Line 215   Column 9   Coefficient -0.02443695
         when "110101101001" => A <= "001001000110101001"; -- Line 215   Column 10   Coefficient 0.14224625
         when "110101101010" => A <= "001000110101000000"; -- Line 215   Column 11   Coefficient 0.13793945
         when "110101101011" => A <= "111111100111100010"; -- Line 215   Column 12   Coefficient -0.00597382
         when "110101101100" => A <= "000000000010010011"; -- Line 215   Column 13   Coefficient 0.00056076
         when "110101101101" => A <= "000000000000000011"; -- Line 215   Column 14   Coefficient 0.00001144
         when "110101101110" => A <= "000000000000000000"; -- Line 215   Column 15   Coefficient 0.00000000
         when "110101101111" => A <= "000000000000000000"; -- Line 215   Column 16   Coefficient 0.00000000
         when "110101110000" => A <= "000000000000000000"; -- Line 216   Column 1   Coefficient 0.00000000
         when "110101110001" => A <= "000000000000000000"; -- Line 216   Column 2   Coefficient 0.00000000
         when "110101110010" => A <= "000000000000000000"; -- Line 216   Column 3   Coefficient 0.00000000
         when "110101110011" => A <= "000000000000000000"; -- Line 216   Column 4   Coefficient 0.00000000
         when "110101110100" => A <= "000000000000000000"; -- Line 216   Column 5   Coefficient 0.00000000
         when "110101110101" => A <= "000000000000000000"; -- Line 216   Column 6   Coefficient 0.00000000
         when "110101110110" => A <= "000000000000000000"; -- Line 216   Column 7   Coefficient 0.00000000
         when "110101110111" => A <= "111111111111001011"; -- Line 216   Column 8   Coefficient -0.00020218
         when "110101111000" => A <= "111110100110010011"; -- Line 216   Column 9   Coefficient -0.02190018
         when "110101111001" => A <= "000111100110110001"; -- Line 216   Column 10   Coefficient 0.11883926
         when "110101111010" => A <= "001010011001111000"; -- Line 216   Column 11   Coefficient 0.16256714
         when "110101111011" => A <= "111111010000101110"; -- Line 216   Column 12   Coefficient -0.01154327
         when "110101111100" => A <= "000000001001011000"; -- Line 216   Column 13   Coefficient 0.00228882
         when "110101111101" => A <= "111111111111110100"; -- Line 216   Column 14   Coefficient -0.00004578
         when "110101111110" => A <= "000000000000000000"; -- Line 216   Column 15   Coefficient 0.00000000
         when "110101111111" => A <= "000000000000000000"; -- Line 216   Column 16   Coefficient 0.00000000
         when "110110000000" => A <= "000000000000000000"; -- Line 217   Column 1   Coefficient 0.00000000
         when "110110000001" => A <= "000000000000000000"; -- Line 217   Column 2   Coefficient 0.00000000
         when "110110000010" => A <= "000000000000000000"; -- Line 217   Column 3   Coefficient 0.00000000
         when "110110000011" => A <= "000000000000000000"; -- Line 217   Column 4   Coefficient 0.00000000
         when "110110000100" => A <= "000000000000000000"; -- Line 217   Column 5   Coefficient 0.00000000
         when "110110000101" => A <= "000000000000000000"; -- Line 217   Column 6   Coefficient 0.00000000
         when "110110000110" => A <= "000000000000000000"; -- Line 217   Column 7   Coefficient 0.00000000
         when "110110000111" => A <= "000000000000000011"; -- Line 217   Column 8   Coefficient 0.00001144
         when "110110001000" => A <= "111110110001100001"; -- Line 217   Column 9   Coefficient -0.01916122
         when "110110001001" => A <= "000110000101110011"; -- Line 217   Column 10   Coefficient 0.09516525
         when "110110001010" => A <= "001011111101111010"; -- Line 217   Column 11   Coefficient 0.18698883
         when "110110001011" => A <= "111110111010000001"; -- Line 217   Column 12   Coefficient -0.01708603
         when "110110001100" => A <= "000000010001001000"; -- Line 217   Column 13   Coefficient 0.00418091
         when "110110001101" => A <= "111111111111100110"; -- Line 217   Column 14   Coefficient -0.00009918
         when "110110001110" => A <= "000000000000000000"; -- Line 217   Column 15   Coefficient 0.00000000
         when "110110001111" => A <= "000000000000000000"; -- Line 217   Column 16   Coefficient 0.00000000
         when "110110010000" => A <= "000000000000000000"; -- Line 218   Column 1   Coefficient 0.00000000
         when "110110010001" => A <= "000000000000000000"; -- Line 218   Column 2   Coefficient 0.00000000
         when "110110010010" => A <= "000000000000000000"; -- Line 218   Column 3   Coefficient 0.00000000
         when "110110010011" => A <= "000000000000000000"; -- Line 218   Column 4   Coefficient 0.00000000
         when "110110010100" => A <= "000000000000000000"; -- Line 218   Column 5   Coefficient 0.00000000
         when "110110010101" => A <= "000000000000000000"; -- Line 218   Column 6   Coefficient 0.00000000
         when "110110010110" => A <= "000000000000000000"; -- Line 218   Column 7   Coefficient 0.00000000
         when "110110010111" => A <= "000000000000001001"; -- Line 218   Column 8   Coefficient 0.00003433
         when "110110011000" => A <= "111111000100111001"; -- Line 218   Column 9   Coefficient -0.01443100
         when "110110011001" => A <= "000100010010000101"; -- Line 218   Column 10   Coefficient 0.06691360
         when "110110011010" => A <= "001101110100101001"; -- Line 218   Column 11   Coefficient 0.21597672
         when "110110011011" => A <= "111110011010010101"; -- Line 218   Column 12   Coefficient -0.02482224
         when "110110011100" => A <= "000000011001110100"; -- Line 218   Column 13   Coefficient 0.00630188
         when "110110011101" => A <= "000000000000000111"; -- Line 218   Column 14   Coefficient 0.00002670
         when "110110011110" => A <= "000000000000000000"; -- Line 218   Column 15   Coefficient 0.00000000
         when "110110011111" => A <= "000000000000000000"; -- Line 218   Column 16   Coefficient 0.00000000
         when "110110100000" => A <= "000000000000000000"; -- Line 219   Column 1   Coefficient 0.00000000
         when "110110100001" => A <= "000000000000000000"; -- Line 219   Column 2   Coefficient 0.00000000
         when "110110100010" => A <= "000000000000000000"; -- Line 219   Column 3   Coefficient 0.00000000
         when "110110100011" => A <= "000000000000000000"; -- Line 219   Column 4   Coefficient 0.00000000
         when "110110100100" => A <= "000000000000000000"; -- Line 219   Column 5   Coefficient 0.00000000
         when "110110100101" => A <= "000000000000000000"; -- Line 219   Column 6   Coefficient 0.00000000
         when "110110100110" => A <= "000000000000000000"; -- Line 219   Column 7   Coefficient 0.00000000
         when "110110100111" => A <= "000000000000000000"; -- Line 219   Column 8   Coefficient 0.00000000
         when "110110101000" => A <= "111111011001111001"; -- Line 219   Column 9   Coefficient -0.00930405
         when "110110101001" => A <= "000010011110111100"; -- Line 219   Column 10   Coefficient 0.03880310
         when "110110101010" => A <= "001111100101110011"; -- Line 219   Column 11   Coefficient 0.24360275
         when "110110101011" => A <= "111101111110110001"; -- Line 219   Column 12   Coefficient -0.03155136
         when "110110101100" => A <= "000000100001110011"; -- Line 219   Column 13   Coefficient 0.00825119
         when "110110101101" => A <= "000000000000110011"; -- Line 219   Column 14   Coefficient 0.00019455
         when "110110101110" => A <= "000000000000000000"; -- Line 219   Column 15   Coefficient 0.00000000
         when "110110101111" => A <= "000000000000000000"; -- Line 219   Column 16   Coefficient 0.00000000
         when "110110110000" => A <= "000000000000000000"; -- Line 220   Column 1   Coefficient 0.00000000
         when "110110110001" => A <= "000000000000000000"; -- Line 220   Column 2   Coefficient 0.00000000
         when "110110110010" => A <= "000000000000000000"; -- Line 220   Column 3   Coefficient 0.00000000
         when "110110110011" => A <= "000000000000000000"; -- Line 220   Column 4   Coefficient 0.00000000
         when "110110110100" => A <= "000000000000000000"; -- Line 220   Column 5   Coefficient 0.00000000
         when "110110110101" => A <= "000000000000000000"; -- Line 220   Column 6   Coefficient 0.00000000
         when "110110110110" => A <= "000000000000000000"; -- Line 220   Column 7   Coefficient 0.00000000
         when "110110110111" => A <= "000000000000000000"; -- Line 220   Column 8   Coefficient 0.00000000
         when "110110111000" => A <= "111111110001010101"; -- Line 220   Column 9   Coefficient -0.00358200
         when "110110111001" => A <= "000000100101011001"; -- Line 220   Column 10   Coefficient 0.00912857
         when "110110111010" => A <= "010001011110001011"; -- Line 220   Column 11   Coefficient 0.27299118
         when "110110111011" => A <= "111101011101101101"; -- Line 220   Column 12   Coefficient -0.03962326
         when "110110111100" => A <= "000000101011110101"; -- Line 220   Column 13   Coefficient 0.01070023
         when "110110111101" => A <= "000000000001100101"; -- Line 220   Column 14   Coefficient 0.00038528
         when "110110111110" => A <= "000000000000000000"; -- Line 220   Column 15   Coefficient 0.00000000
         when "110110111111" => A <= "000000000000000000"; -- Line 220   Column 16   Coefficient 0.00000000
         when "110111000000" => A <= "000000000000000000"; -- Line 221   Column 1   Coefficient 0.00000000
         when "110111000001" => A <= "000000000000000000"; -- Line 221   Column 2   Coefficient 0.00000000
         when "110111000010" => A <= "000000000000000000"; -- Line 221   Column 3   Coefficient 0.00000000
         when "110111000011" => A <= "000000000000000000"; -- Line 221   Column 4   Coefficient 0.00000000
         when "110111000100" => A <= "000000000000000000"; -- Line 221   Column 5   Coefficient 0.00000000
         when "110111000101" => A <= "000000000000000000"; -- Line 221   Column 6   Coefficient 0.00000000
         when "110111000110" => A <= "000000000000000000"; -- Line 221   Column 7   Coefficient 0.00000000
         when "110111000111" => A <= "000000000000000000"; -- Line 221   Column 8   Coefficient 0.00000000
         when "110111001000" => A <= "000000000111011010"; -- Line 221   Column 9   Coefficient 0.00180817
         when "110111001001" => A <= "111110110101100100"; -- Line 221   Column 10   Coefficient -0.01817322
         when "110111001010" => A <= "010011000101100111"; -- Line 221   Column 11   Coefficient 0.29824448
         when "110111001011" => A <= "111101000110110001"; -- Line 221   Column 12   Coefficient -0.04522324
         when "110111001100" => A <= "000000110100010110"; -- Line 221   Column 13   Coefficient 0.01277924
         when "110111001101" => A <= "000000000010010101"; -- Line 221   Column 14   Coefficient 0.00056839
         when "110111001110" => A <= "000000000000000000"; -- Line 221   Column 15   Coefficient 0.00000000
         when "110111001111" => A <= "000000000000000000"; -- Line 221   Column 16   Coefficient 0.00000000
         when "110111010000" => A <= "000000000000000000"; -- Line 222   Column 1   Coefficient 0.00000000
         when "110111010001" => A <= "000000000000000000"; -- Line 222   Column 2   Coefficient 0.00000000
         when "110111010010" => A <= "000000000000000000"; -- Line 222   Column 3   Coefficient 0.00000000
         when "110111010011" => A <= "000000000000000000"; -- Line 222   Column 4   Coefficient 0.00000000
         when "110111010100" => A <= "000000000000000000"; -- Line 222   Column 5   Coefficient 0.00000000
         when "110111010101" => A <= "000000000000000000"; -- Line 222   Column 6   Coefficient 0.00000000
         when "110111010110" => A <= "000000000000000000"; -- Line 222   Column 7   Coefficient 0.00000000
         when "110111010111" => A <= "000000000000000000"; -- Line 222   Column 8   Coefficient 0.00000000
         when "110111011000" => A <= "000000001111000010"; -- Line 222   Column 9   Coefficient 0.00366974
         when "110111011001" => A <= "111110000010011110"; -- Line 222   Column 10   Coefficient -0.03064728
         when "110111011010" => A <= "010011010010100110"; -- Line 222   Column 11   Coefficient 0.30141449
         when "110111011011" => A <= "111101100111001110"; -- Line 222   Column 12   Coefficient -0.03730011
         when "110111011100" => A <= "000000110010101110"; -- Line 222   Column 13   Coefficient 0.01238251
         when "110111011101" => A <= "000000000001111110"; -- Line 222   Column 14   Coefficient 0.00048065
         when "110111011110" => A <= "000000000000000000"; -- Line 222   Column 15   Coefficient 0.00000000
         when "110111011111" => A <= "000000000000000000"; -- Line 222   Column 16   Coefficient 0.00000000
         when "110111100000" => A <= "000000000000000000"; -- Line 223   Column 1   Coefficient 0.00000000
         when "110111100001" => A <= "000000000000000000"; -- Line 223   Column 2   Coefficient 0.00000000
         when "110111100010" => A <= "000000000000000000"; -- Line 223   Column 3   Coefficient 0.00000000
         when "110111100011" => A <= "000000000000000000"; -- Line 223   Column 4   Coefficient 0.00000000
         when "110111100100" => A <= "000000000000000000"; -- Line 223   Column 5   Coefficient 0.00000000
         when "110111100101" => A <= "000000000000000000"; -- Line 223   Column 6   Coefficient 0.00000000
         when "110111100110" => A <= "000000000000000000"; -- Line 223   Column 7   Coefficient 0.00000000
         when "110111100111" => A <= "000000000000000000"; -- Line 223   Column 8   Coefficient 0.00000000
         when "110111101000" => A <= "000000010000011000"; -- Line 223   Column 9   Coefficient 0.00399780
         when "110111101001" => A <= "111101101011101110"; -- Line 223   Column 10   Coefficient -0.03620148
         when "110111101010" => A <= "010010110100110100"; -- Line 223   Column 11   Coefficient 0.29414368
         when "110111101011" => A <= "111110100000101100"; -- Line 223   Column 12   Coefficient -0.02326965
         when "110111101100" => A <= "000000101101010111"; -- Line 223   Column 13   Coefficient 0.01107407
         when "110111101101" => A <= "000000000001000010"; -- Line 223   Column 14   Coefficient 0.00025177
         when "110111101110" => A <= "000000000000000000"; -- Line 223   Column 15   Coefficient 0.00000000
         when "110111101111" => A <= "000000000000000000"; -- Line 223   Column 16   Coefficient 0.00000000
         when "110111110000" => A <= "000000000000000000"; -- Line 224   Column 1   Coefficient 0.00000000
         when "110111110001" => A <= "000000000000000000"; -- Line 224   Column 2   Coefficient 0.00000000
         when "110111110010" => A <= "000000000000000000"; -- Line 224   Column 3   Coefficient 0.00000000
         when "110111110011" => A <= "000000000000000000"; -- Line 224   Column 4   Coefficient 0.00000000
         when "110111110100" => A <= "000000000000000000"; -- Line 224   Column 5   Coefficient 0.00000000
         when "110111110101" => A <= "000000000000000000"; -- Line 224   Column 6   Coefficient 0.00000000
         when "110111110110" => A <= "000000000000000000"; -- Line 224   Column 7   Coefficient 0.00000000
         when "110111110111" => A <= "000000000000000000"; -- Line 224   Column 8   Coefficient 0.00000000
         when "110111111000" => A <= "000000001111111100"; -- Line 224   Column 9   Coefficient 0.00389099
         when "110111111001" => A <= "111101100000101101"; -- Line 224   Column 10   Coefficient -0.03889084
         when "110111111010" => A <= "010010000001100011"; -- Line 224   Column 11   Coefficient 0.28162766
         when "110111111011" => A <= "111111101010001000"; -- Line 224   Column 12   Coefficient -0.00534058
         when "110111111100" => A <= "000000100010100100"; -- Line 224   Column 13   Coefficient 0.00843811
         when "110111111101" => A <= "000000000001001000"; -- Line 224   Column 14   Coefficient 0.00027466
         when "110111111110" => A <= "000000000000000000"; -- Line 224   Column 15   Coefficient 0.00000000
         when "110111111111" => A <= "000000000000000000"; -- Line 224   Column 16   Coefficient 0.00000000
         when "111000000000" => A <= "000000000000000000"; -- Line 225   Column 1   Coefficient 0.00000000
         when "111000000001" => A <= "000000000000000000"; -- Line 225   Column 2   Coefficient 0.00000000
         when "111000000010" => A <= "000000000000000000"; -- Line 225   Column 3   Coefficient 0.00000000
         when "111000000011" => A <= "000000000000000000"; -- Line 225   Column 4   Coefficient 0.00000000
         when "111000000100" => A <= "000000000000000000"; -- Line 225   Column 5   Coefficient 0.00000000
         when "111000000101" => A <= "000000000000000000"; -- Line 225   Column 6   Coefficient 0.00000000
         when "111000000110" => A <= "000000000000000000"; -- Line 225   Column 7   Coefficient 0.00000000
         when "111000000111" => A <= "000000000000000000"; -- Line 225   Column 8   Coefficient 0.00000000
         when "111000001000" => A <= "000000001101001100"; -- Line 225   Column 9   Coefficient 0.00321960
         when "111000001001" => A <= "111101100010001110"; -- Line 225   Column 10   Coefficient -0.03852081
         when "111000001010" => A <= "010000111010100101"; -- Line 225   Column 11   Coefficient 0.26430130
         when "111000001011" => A <= "000000111110100110"; -- Line 225   Column 12   Coefficient 0.01528168
         when "111000001100" => A <= "000000010110010000"; -- Line 225   Column 13   Coefficient 0.00543213
         when "111000001101" => A <= "000000000001001011"; -- Line 225   Column 14   Coefficient 0.00028610
         when "111000001110" => A <= "000000000000000000"; -- Line 225   Column 15   Coefficient 0.00000000
         when "111000001111" => A <= "000000000000000000"; -- Line 225   Column 16   Coefficient 0.00000000
         when "111000010000" => A <= "000000000000000000"; -- Line 226   Column 1   Coefficient 0.00000000
         when "111000010001" => A <= "000000000000000000"; -- Line 226   Column 2   Coefficient 0.00000000
         when "111000010010" => A <= "000000000000000000"; -- Line 226   Column 3   Coefficient 0.00000000
         when "111000010011" => A <= "000000000000000000"; -- Line 226   Column 4   Coefficient 0.00000000
         when "111000010100" => A <= "000000000000000000"; -- Line 226   Column 5   Coefficient 0.00000000
         when "111000010101" => A <= "000000000000000000"; -- Line 226   Column 6   Coefficient 0.00000000
         when "111000010110" => A <= "000000000000000000"; -- Line 226   Column 7   Coefficient 0.00000000
         when "111000010111" => A <= "000000000000000000"; -- Line 226   Column 8   Coefficient 0.00000000
         when "111000011000" => A <= "000000001010110110"; -- Line 226   Column 9   Coefficient 0.00264740
         when "111000011001" => A <= "111101100010101111"; -- Line 226   Column 10   Coefficient -0.03839493
         when "111000011010" => A <= "001111111010100001"; -- Line 226   Column 11   Coefficient 0.24866104
         when "111000011011" => A <= "000010000100001011"; -- Line 226   Column 12   Coefficient 0.03226852
         when "111000011100" => A <= "000000010100110111"; -- Line 226   Column 13   Coefficient 0.00509262
         when "111000011101" => A <= "111111111110110111"; -- Line 226   Column 14   Coefficient -0.00027847
         when "111000011110" => A <= "000000000000000000"; -- Line 226   Column 15   Coefficient 0.00000000
         when "111000011111" => A <= "000000000000000000"; -- Line 226   Column 16   Coefficient 0.00000000
         when "111000100000" => A <= "000000000000000000"; -- Line 227   Column 1   Coefficient 0.00000000
         when "111000100001" => A <= "000000000000000000"; -- Line 227   Column 2   Coefficient 0.00000000
         when "111000100010" => A <= "000000000000000000"; -- Line 227   Column 3   Coefficient 0.00000000
         when "111000100011" => A <= "000000000000000000"; -- Line 227   Column 4   Coefficient 0.00000000
         when "111000100100" => A <= "000000000000000000"; -- Line 227   Column 5   Coefficient 0.00000000
         when "111000100101" => A <= "000000000000000000"; -- Line 227   Column 6   Coefficient 0.00000000
         when "111000100110" => A <= "000000000000000000"; -- Line 227   Column 7   Coefficient 0.00000000
         when "111000100111" => A <= "000000000000000000"; -- Line 227   Column 8   Coefficient 0.00000000
         when "111000101000" => A <= "000000001000010011"; -- Line 227   Column 9   Coefficient 0.00202560
         when "111000101001" => A <= "111101100110110000"; -- Line 227   Column 10   Coefficient -0.03741455
         when "111000101010" => A <= "001110110101010100"; -- Line 227   Column 11   Coefficient 0.23176575
         when "111000101011" => A <= "000011001010010011"; -- Line 227   Column 12   Coefficient 0.04938889
         when "111000101100" => A <= "000000010100111001"; -- Line 227   Column 13   Coefficient 0.00510025
         when "111000101101" => A <= "111111111100011110"; -- Line 227   Column 14   Coefficient -0.00086212
         when "111000101110" => A <= "111111111111111111"; -- Line 227   Column 15   Coefficient -0.00000381
         when "111000101111" => A <= "000000000000000000"; -- Line 227   Column 16   Coefficient 0.00000000
         when "111000110000" => A <= "000000000000000000"; -- Line 228   Column 1   Coefficient 0.00000000
         when "111000110001" => A <= "000000000000000000"; -- Line 228   Column 2   Coefficient 0.00000000
         when "111000110010" => A <= "000000000000000000"; -- Line 228   Column 3   Coefficient 0.00000000
         when "111000110011" => A <= "000000000000000000"; -- Line 228   Column 4   Coefficient 0.00000000
         when "111000110100" => A <= "000000000000000000"; -- Line 228   Column 5   Coefficient 0.00000000
         when "111000110101" => A <= "000000000000000000"; -- Line 228   Column 6   Coefficient 0.00000000
         when "111000110110" => A <= "000000000000000000"; -- Line 228   Column 7   Coefficient 0.00000000
         when "111000110111" => A <= "000000000000000000"; -- Line 228   Column 8   Coefficient 0.00000000
         when "111000111000" => A <= "000000000011111000"; -- Line 228   Column 9   Coefficient 0.00094604
         when "111000111001" => A <= "111101110100001010"; -- Line 228   Column 10   Coefficient -0.03414154
         when "111000111010" => A <= "001101100011111111"; -- Line 228   Column 11   Coefficient 0.21191025
         when "111000111011" => A <= "000100010011001101"; -- Line 228   Column 12   Coefficient 0.06718826
         when "111000111100" => A <= "000000010111101010"; -- Line 228   Column 13   Coefficient 0.00577545
         when "111000111101" => A <= "111111111001000110"; -- Line 228   Column 14   Coefficient -0.00168610
         when "111000111110" => A <= "000000000000000011"; -- Line 228   Column 15   Coefficient 0.00001144
         when "111000111111" => A <= "000000000000000000"; -- Line 228   Column 16   Coefficient 0.00000000
         when "111001000000" => A <= "000000000000000000"; -- Line 229   Column 1   Coefficient 0.00000000
         when "111001000001" => A <= "000000000000000000"; -- Line 229   Column 2   Coefficient 0.00000000
         when "111001000010" => A <= "000000000000000000"; -- Line 229   Column 3   Coefficient 0.00000000
         when "111001000011" => A <= "000000000000000000"; -- Line 229   Column 4   Coefficient 0.00000000
         when "111001000100" => A <= "000000000000000000"; -- Line 229   Column 5   Coefficient 0.00000000
         when "111001000101" => A <= "000000000000000000"; -- Line 229   Column 6   Coefficient 0.00000000
         when "111001000110" => A <= "000000000000000000"; -- Line 229   Column 7   Coefficient 0.00000000
         when "111001000111" => A <= "000000000000000000"; -- Line 229   Column 8   Coefficient 0.00000000
         when "111001001000" => A <= "111111111111010011"; -- Line 229   Column 9   Coefficient -0.00017166
         when "111001001001" => A <= "111110000101010011"; -- Line 229   Column 10   Coefficient -0.02995682
         when "111001001010" => A <= "001100001011101000"; -- Line 229   Column 11   Coefficient 0.19033813
         when "111001001011" => A <= "000101100000010101"; -- Line 229   Column 12   Coefficient 0.08601761
         when "111001001100" => A <= "000000011000110111"; -- Line 229   Column 13   Coefficient 0.00606918
         when "111001001101" => A <= "111111110110011111"; -- Line 229   Column 14   Coefficient -0.00232315
         when "111001001110" => A <= "000000000000000110"; -- Line 229   Column 15   Coefficient 0.00002289
         when "111001001111" => A <= "000000000000000000"; -- Line 229   Column 16   Coefficient 0.00000000
         when "111001010000" => A <= "000000000000000000"; -- Line 230   Column 1   Coefficient 0.00000000
         when "111001010001" => A <= "000000000000000000"; -- Line 230   Column 2   Coefficient 0.00000000
         when "111001010010" => A <= "000000000000000000"; -- Line 230   Column 3   Coefficient 0.00000000
         when "111001010011" => A <= "000000000000000000"; -- Line 230   Column 4   Coefficient 0.00000000
         when "111001010100" => A <= "000000000000000000"; -- Line 230   Column 5   Coefficient 0.00000000
         when "111001010101" => A <= "000000000000000000"; -- Line 230   Column 6   Coefficient 0.00000000
         when "111001010110" => A <= "000000000000000000"; -- Line 230   Column 7   Coefficient 0.00000000
         when "111001010111" => A <= "000000000000000000"; -- Line 230   Column 8   Coefficient 0.00000000
         when "111001011000" => A <= "111111111110010010"; -- Line 230   Column 9   Coefficient -0.00041962
         when "111001011001" => A <= "111110010000110000"; -- Line 230   Column 10   Coefficient -0.02716064
         when "111001011010" => A <= "001010101100000111"; -- Line 230   Column 11   Coefficient 0.16701889
         when "111001011011" => A <= "000111000101010101"; -- Line 230   Column 12   Coefficient 0.11067581
         when "111001011100" => A <= "000000000100100100"; -- Line 230   Column 13   Coefficient 0.00111389
         when "111001011101" => A <= "111111111010111001"; -- Line 230   Column 14   Coefficient -0.00124741
         when "111001011110" => A <= "000000000000000100"; -- Line 230   Column 15   Coefficient 0.00001526
         when "111001011111" => A <= "000000000000000000"; -- Line 230   Column 16   Coefficient 0.00000000
         when "111001100000" => A <= "000000000000000000"; -- Line 231   Column 1   Coefficient 0.00000000
         when "111001100001" => A <= "000000000000000000"; -- Line 231   Column 2   Coefficient 0.00000000
         when "111001100010" => A <= "000000000000000000"; -- Line 231   Column 3   Coefficient 0.00000000
         when "111001100011" => A <= "000000000000000000"; -- Line 231   Column 4   Coefficient 0.00000000
         when "111001100100" => A <= "000000000000000000"; -- Line 231   Column 5   Coefficient 0.00000000
         when "111001100101" => A <= "000000000000000000"; -- Line 231   Column 6   Coefficient 0.00000000
         when "111001100110" => A <= "000000000000000000"; -- Line 231   Column 7   Coefficient 0.00000000
         when "111001100111" => A <= "000000000000000000"; -- Line 231   Column 8   Coefficient 0.00000000
         when "111001101000" => A <= "111111111110100110"; -- Line 231   Column 9   Coefficient -0.00034332
         when "111001101001" => A <= "111110011011111010"; -- Line 231   Column 10   Coefficient -0.02443695
         when "111001101010" => A <= "001001000110101001"; -- Line 231   Column 11   Coefficient 0.14224625
         when "111001101011" => A <= "001000110101000000"; -- Line 231   Column 12   Coefficient 0.13793945
         when "111001101100" => A <= "111111100111100010"; -- Line 231   Column 13   Coefficient -0.00597382
         when "111001101101" => A <= "000000000010010011"; -- Line 231   Column 14   Coefficient 0.00056076
         when "111001101110" => A <= "000000000000000011"; -- Line 231   Column 15   Coefficient 0.00001144
         when "111001101111" => A <= "000000000000000000"; -- Line 231   Column 16   Coefficient 0.00000000
         when "111001110000" => A <= "000000000000000000"; -- Line 232   Column 1   Coefficient 0.00000000
         when "111001110001" => A <= "000000000000000000"; -- Line 232   Column 2   Coefficient 0.00000000
         when "111001110010" => A <= "000000000000000000"; -- Line 232   Column 3   Coefficient 0.00000000
         when "111001110011" => A <= "000000000000000000"; -- Line 232   Column 4   Coefficient 0.00000000
         when "111001110100" => A <= "000000000000000000"; -- Line 232   Column 5   Coefficient 0.00000000
         when "111001110101" => A <= "000000000000000000"; -- Line 232   Column 6   Coefficient 0.00000000
         when "111001110110" => A <= "000000000000000000"; -- Line 232   Column 7   Coefficient 0.00000000
         when "111001110111" => A <= "000000000000000000"; -- Line 232   Column 8   Coefficient 0.00000000
         when "111001111000" => A <= "111111111111001011"; -- Line 232   Column 9   Coefficient -0.00020218
         when "111001111001" => A <= "111110100110010011"; -- Line 232   Column 10   Coefficient -0.02190018
         when "111001111010" => A <= "000111100110110001"; -- Line 232   Column 11   Coefficient 0.11883926
         when "111001111011" => A <= "001010011001111000"; -- Line 232   Column 12   Coefficient 0.16256714
         when "111001111100" => A <= "111111010000101110"; -- Line 232   Column 13   Coefficient -0.01154327
         when "111001111101" => A <= "000000001001011000"; -- Line 232   Column 14   Coefficient 0.00228882
         when "111001111110" => A <= "111111111111110100"; -- Line 232   Column 15   Coefficient -0.00004578
         when "111001111111" => A <= "000000000000000000"; -- Line 232   Column 16   Coefficient 0.00000000
         when "111010000000" => A <= "000000000000000000"; -- Line 233   Column 1   Coefficient 0.00000000
         when "111010000001" => A <= "000000000000000000"; -- Line 233   Column 2   Coefficient 0.00000000
         when "111010000010" => A <= "000000000000000000"; -- Line 233   Column 3   Coefficient 0.00000000
         when "111010000011" => A <= "000000000000000000"; -- Line 233   Column 4   Coefficient 0.00000000
         when "111010000100" => A <= "000000000000000000"; -- Line 233   Column 5   Coefficient 0.00000000
         when "111010000101" => A <= "000000000000000000"; -- Line 233   Column 6   Coefficient 0.00000000
         when "111010000110" => A <= "000000000000000000"; -- Line 233   Column 7   Coefficient 0.00000000
         when "111010000111" => A <= "000000000000000000"; -- Line 233   Column 8   Coefficient 0.00000000
         when "111010001000" => A <= "000000000000000011"; -- Line 233   Column 9   Coefficient 0.00001144
         when "111010001001" => A <= "111110110001100001"; -- Line 233   Column 10   Coefficient -0.01916122
         when "111010001010" => A <= "000110000101110011"; -- Line 233   Column 11   Coefficient 0.09516525
         when "111010001011" => A <= "001011111101111010"; -- Line 233   Column 12   Coefficient 0.18698883
         when "111010001100" => A <= "111110111010000001"; -- Line 233   Column 13   Coefficient -0.01708603
         when "111010001101" => A <= "000000010001001000"; -- Line 233   Column 14   Coefficient 0.00418091
         when "111010001110" => A <= "111111111111100110"; -- Line 233   Column 15   Coefficient -0.00009918
         when "111010001111" => A <= "000000000000000000"; -- Line 233   Column 16   Coefficient 0.00000000
         when "111010010000" => A <= "000000000000000000"; -- Line 234   Column 1   Coefficient 0.00000000
         when "111010010001" => A <= "000000000000000000"; -- Line 234   Column 2   Coefficient 0.00000000
         when "111010010010" => A <= "000000000000000000"; -- Line 234   Column 3   Coefficient 0.00000000
         when "111010010011" => A <= "000000000000000000"; -- Line 234   Column 4   Coefficient 0.00000000
         when "111010010100" => A <= "000000000000000000"; -- Line 234   Column 5   Coefficient 0.00000000
         when "111010010101" => A <= "000000000000000000"; -- Line 234   Column 6   Coefficient 0.00000000
         when "111010010110" => A <= "000000000000000000"; -- Line 234   Column 7   Coefficient 0.00000000
         when "111010010111" => A <= "000000000000000000"; -- Line 234   Column 8   Coefficient 0.00000000
         when "111010011000" => A <= "000000000000001001"; -- Line 234   Column 9   Coefficient 0.00003433
         when "111010011001" => A <= "111111000100111001"; -- Line 234   Column 10   Coefficient -0.01443100
         when "111010011010" => A <= "000100010010000101"; -- Line 234   Column 11   Coefficient 0.06691360
         when "111010011011" => A <= "001101110100101001"; -- Line 234   Column 12   Coefficient 0.21597672
         when "111010011100" => A <= "111110011010010101"; -- Line 234   Column 13   Coefficient -0.02482224
         when "111010011101" => A <= "000000011001110100"; -- Line 234   Column 14   Coefficient 0.00630188
         when "111010011110" => A <= "000000000000000111"; -- Line 234   Column 15   Coefficient 0.00002670
         when "111010011111" => A <= "000000000000000000"; -- Line 234   Column 16   Coefficient 0.00000000
         when "111010100000" => A <= "000000000000000000"; -- Line 235   Column 1   Coefficient 0.00000000
         when "111010100001" => A <= "000000000000000000"; -- Line 235   Column 2   Coefficient 0.00000000
         when "111010100010" => A <= "000000000000000000"; -- Line 235   Column 3   Coefficient 0.00000000
         when "111010100011" => A <= "000000000000000000"; -- Line 235   Column 4   Coefficient 0.00000000
         when "111010100100" => A <= "000000000000000000"; -- Line 235   Column 5   Coefficient 0.00000000
         when "111010100101" => A <= "000000000000000000"; -- Line 235   Column 6   Coefficient 0.00000000
         when "111010100110" => A <= "000000000000000000"; -- Line 235   Column 7   Coefficient 0.00000000
         when "111010100111" => A <= "000000000000000000"; -- Line 235   Column 8   Coefficient 0.00000000
         when "111010101000" => A <= "000000000000000000"; -- Line 235   Column 9   Coefficient 0.00000000
         when "111010101001" => A <= "111111011001111001"; -- Line 235   Column 10   Coefficient -0.00930405
         when "111010101010" => A <= "000010011110111100"; -- Line 235   Column 11   Coefficient 0.03880310
         when "111010101011" => A <= "001111100101110011"; -- Line 235   Column 12   Coefficient 0.24360275
         when "111010101100" => A <= "111101111110110001"; -- Line 235   Column 13   Coefficient -0.03155136
         when "111010101101" => A <= "000000100001110011"; -- Line 235   Column 14   Coefficient 0.00825119
         when "111010101110" => A <= "000000000000110011"; -- Line 235   Column 15   Coefficient 0.00019455
         when "111010101111" => A <= "000000000000000000"; -- Line 235   Column 16   Coefficient 0.00000000
         when "111010110000" => A <= "000000000000000000"; -- Line 236   Column 1   Coefficient 0.00000000
         when "111010110001" => A <= "000000000000000000"; -- Line 236   Column 2   Coefficient 0.00000000
         when "111010110010" => A <= "000000000000000000"; -- Line 236   Column 3   Coefficient 0.00000000
         when "111010110011" => A <= "000000000000000000"; -- Line 236   Column 4   Coefficient 0.00000000
         when "111010110100" => A <= "000000000000000000"; -- Line 236   Column 5   Coefficient 0.00000000
         when "111010110101" => A <= "000000000000000000"; -- Line 236   Column 6   Coefficient 0.00000000
         when "111010110110" => A <= "000000000000000000"; -- Line 236   Column 7   Coefficient 0.00000000
         when "111010110111" => A <= "000000000000000000"; -- Line 236   Column 8   Coefficient 0.00000000
         when "111010111000" => A <= "000000000000000000"; -- Line 236   Column 9   Coefficient 0.00000000
         when "111010111001" => A <= "111111110001010101"; -- Line 236   Column 10   Coefficient -0.00358200
         when "111010111010" => A <= "000000100101011001"; -- Line 236   Column 11   Coefficient 0.00912857
         when "111010111011" => A <= "010001011110001011"; -- Line 236   Column 12   Coefficient 0.27299118
         when "111010111100" => A <= "111101011101101101"; -- Line 236   Column 13   Coefficient -0.03962326
         when "111010111101" => A <= "000000101011110101"; -- Line 236   Column 14   Coefficient 0.01070023
         when "111010111110" => A <= "000000000001100101"; -- Line 236   Column 15   Coefficient 0.00038528
         when "111010111111" => A <= "000000000000000000"; -- Line 236   Column 16   Coefficient 0.00000000
         when "111011000000" => A <= "000000000000000000"; -- Line 237   Column 1   Coefficient 0.00000000
         when "111011000001" => A <= "000000000000000000"; -- Line 237   Column 2   Coefficient 0.00000000
         when "111011000010" => A <= "000000000000000000"; -- Line 237   Column 3   Coefficient 0.00000000
         when "111011000011" => A <= "000000000000000000"; -- Line 237   Column 4   Coefficient 0.00000000
         when "111011000100" => A <= "000000000000000000"; -- Line 237   Column 5   Coefficient 0.00000000
         when "111011000101" => A <= "000000000000000000"; -- Line 237   Column 6   Coefficient 0.00000000
         when "111011000110" => A <= "000000000000000000"; -- Line 237   Column 7   Coefficient 0.00000000
         when "111011000111" => A <= "000000000000000000"; -- Line 237   Column 8   Coefficient 0.00000000
         when "111011001000" => A <= "000000000000000000"; -- Line 237   Column 9   Coefficient 0.00000000
         when "111011001001" => A <= "000000000111011010"; -- Line 237   Column 10   Coefficient 0.00180817
         when "111011001010" => A <= "111110110101100100"; -- Line 237   Column 11   Coefficient -0.01817322
         when "111011001011" => A <= "010011000101100111"; -- Line 237   Column 12   Coefficient 0.29824448
         when "111011001100" => A <= "111101000110110001"; -- Line 237   Column 13   Coefficient -0.04522324
         when "111011001101" => A <= "000000110100010110"; -- Line 237   Column 14   Coefficient 0.01277924
         when "111011001110" => A <= "000000000010010101"; -- Line 237   Column 15   Coefficient 0.00056839
         when "111011001111" => A <= "000000000000000000"; -- Line 237   Column 16   Coefficient 0.00000000
         when "111011010000" => A <= "000000000000000000"; -- Line 238   Column 1   Coefficient 0.00000000
         when "111011010001" => A <= "000000000000000000"; -- Line 238   Column 2   Coefficient 0.00000000
         when "111011010010" => A <= "000000000000000000"; -- Line 238   Column 3   Coefficient 0.00000000
         when "111011010011" => A <= "000000000000000000"; -- Line 238   Column 4   Coefficient 0.00000000
         when "111011010100" => A <= "000000000000000000"; -- Line 238   Column 5   Coefficient 0.00000000
         when "111011010101" => A <= "000000000000000000"; -- Line 238   Column 6   Coefficient 0.00000000
         when "111011010110" => A <= "000000000000000000"; -- Line 238   Column 7   Coefficient 0.00000000
         when "111011010111" => A <= "000000000000000000"; -- Line 238   Column 8   Coefficient 0.00000000
         when "111011011000" => A <= "000000000000000000"; -- Line 238   Column 9   Coefficient 0.00000000
         when "111011011001" => A <= "000000001111000010"; -- Line 238   Column 10   Coefficient 0.00366974
         when "111011011010" => A <= "111110000010011110"; -- Line 238   Column 11   Coefficient -0.03064728
         when "111011011011" => A <= "010011010010100110"; -- Line 238   Column 12   Coefficient 0.30141449
         when "111011011100" => A <= "111101100111001110"; -- Line 238   Column 13   Coefficient -0.03730011
         when "111011011101" => A <= "000000110010101110"; -- Line 238   Column 14   Coefficient 0.01238251
         when "111011011110" => A <= "000000000001111110"; -- Line 238   Column 15   Coefficient 0.00048065
         when "111011011111" => A <= "000000000000000000"; -- Line 238   Column 16   Coefficient 0.00000000
         when "111011100000" => A <= "000000000000000000"; -- Line 239   Column 1   Coefficient 0.00000000
         when "111011100001" => A <= "000000000000000000"; -- Line 239   Column 2   Coefficient 0.00000000
         when "111011100010" => A <= "000000000000000000"; -- Line 239   Column 3   Coefficient 0.00000000
         when "111011100011" => A <= "000000000000000000"; -- Line 239   Column 4   Coefficient 0.00000000
         when "111011100100" => A <= "000000000000000000"; -- Line 239   Column 5   Coefficient 0.00000000
         when "111011100101" => A <= "000000000000000000"; -- Line 239   Column 6   Coefficient 0.00000000
         when "111011100110" => A <= "000000000000000000"; -- Line 239   Column 7   Coefficient 0.00000000
         when "111011100111" => A <= "000000000000000000"; -- Line 239   Column 8   Coefficient 0.00000000
         when "111011101000" => A <= "000000000000000000"; -- Line 239   Column 9   Coefficient 0.00000000
         when "111011101001" => A <= "000000010000011000"; -- Line 239   Column 10   Coefficient 0.00399780
         when "111011101010" => A <= "111101101011101110"; -- Line 239   Column 11   Coefficient -0.03620148
         when "111011101011" => A <= "010010110100110100"; -- Line 239   Column 12   Coefficient 0.29414368
         when "111011101100" => A <= "111110100000101100"; -- Line 239   Column 13   Coefficient -0.02326965
         when "111011101101" => A <= "000000101101010111"; -- Line 239   Column 14   Coefficient 0.01107407
         when "111011101110" => A <= "000000000001000010"; -- Line 239   Column 15   Coefficient 0.00025177
         when "111011101111" => A <= "000000000000000000"; -- Line 239   Column 16   Coefficient 0.00000000
         when "111011110000" => A <= "000000000000000000"; -- Line 240   Column 1   Coefficient 0.00000000
         when "111011110001" => A <= "000000000000000000"; -- Line 240   Column 2   Coefficient 0.00000000
         when "111011110010" => A <= "000000000000000000"; -- Line 240   Column 3   Coefficient 0.00000000
         when "111011110011" => A <= "000000000000000000"; -- Line 240   Column 4   Coefficient 0.00000000
         when "111011110100" => A <= "000000000000000000"; -- Line 240   Column 5   Coefficient 0.00000000
         when "111011110101" => A <= "000000000000000000"; -- Line 240   Column 6   Coefficient 0.00000000
         when "111011110110" => A <= "000000000000000000"; -- Line 240   Column 7   Coefficient 0.00000000
         when "111011110111" => A <= "000000000000000000"; -- Line 240   Column 8   Coefficient 0.00000000
         when "111011111000" => A <= "000000000000000000"; -- Line 240   Column 9   Coefficient 0.00000000
         when "111011111001" => A <= "000000001111111100"; -- Line 240   Column 10   Coefficient 0.00389099
         when "111011111010" => A <= "111101100000101101"; -- Line 240   Column 11   Coefficient -0.03889084
         when "111011111011" => A <= "010010000001100011"; -- Line 240   Column 12   Coefficient 0.28162766
         when "111011111100" => A <= "111111101010001000"; -- Line 240   Column 13   Coefficient -0.00534058
         when "111011111101" => A <= "000000100010100100"; -- Line 240   Column 14   Coefficient 0.00843811
         when "111011111110" => A <= "000000000001001000"; -- Line 240   Column 15   Coefficient 0.00027466
         when "111011111111" => A <= "000000000000000000"; -- Line 240   Column 16   Coefficient 0.00000000
         when "111100000000" => A <= "000000000000000000"; -- Line 241   Column 1   Coefficient 0.00000000
         when "111100000001" => A <= "000000000000000000"; -- Line 241   Column 2   Coefficient 0.00000000
         when "111100000010" => A <= "000000000000000000"; -- Line 241   Column 3   Coefficient 0.00000000
         when "111100000011" => A <= "000000000000000000"; -- Line 241   Column 4   Coefficient 0.00000000
         when "111100000100" => A <= "000000000000000000"; -- Line 241   Column 5   Coefficient 0.00000000
         when "111100000101" => A <= "000000000000000000"; -- Line 241   Column 6   Coefficient 0.00000000
         when "111100000110" => A <= "000000000000000000"; -- Line 241   Column 7   Coefficient 0.00000000
         when "111100000111" => A <= "000000000000000000"; -- Line 241   Column 8   Coefficient 0.00000000
         when "111100001000" => A <= "000000000000000000"; -- Line 241   Column 9   Coefficient 0.00000000
         when "111100001001" => A <= "000000001101001100"; -- Line 241   Column 10   Coefficient 0.00321960
         when "111100001010" => A <= "111101100010001110"; -- Line 241   Column 11   Coefficient -0.03852081
         when "111100001011" => A <= "010000111010100101"; -- Line 241   Column 12   Coefficient 0.26430130
         when "111100001100" => A <= "000000111110100110"; -- Line 241   Column 13   Coefficient 0.01528168
         when "111100001101" => A <= "000000010110010000"; -- Line 241   Column 14   Coefficient 0.00543213
         when "111100001110" => A <= "000000000001001011"; -- Line 241   Column 15   Coefficient 0.00028610
         when "111100001111" => A <= "000000000000000000"; -- Line 241   Column 16   Coefficient 0.00000000
         when "111100010000" => A <= "000000000000000000"; -- Line 242   Column 1   Coefficient 0.00000000
         when "111100010001" => A <= "000000000000000000"; -- Line 242   Column 2   Coefficient 0.00000000
         when "111100010010" => A <= "000000000000000000"; -- Line 242   Column 3   Coefficient 0.00000000
         when "111100010011" => A <= "000000000000000000"; -- Line 242   Column 4   Coefficient 0.00000000
         when "111100010100" => A <= "000000000000000000"; -- Line 242   Column 5   Coefficient 0.00000000
         when "111100010101" => A <= "000000000000000000"; -- Line 242   Column 6   Coefficient 0.00000000
         when "111100010110" => A <= "000000000000000000"; -- Line 242   Column 7   Coefficient 0.00000000
         when "111100010111" => A <= "000000000000000000"; -- Line 242   Column 8   Coefficient 0.00000000
         when "111100011000" => A <= "000000000000000000"; -- Line 242   Column 9   Coefficient 0.00000000
         when "111100011001" => A <= "000000001010110110"; -- Line 242   Column 10   Coefficient 0.00264740
         when "111100011010" => A <= "111101100010101111"; -- Line 242   Column 11   Coefficient -0.03839493
         when "111100011011" => A <= "001111111010100001"; -- Line 242   Column 12   Coefficient 0.24866104
         when "111100011100" => A <= "000010000100001011"; -- Line 242   Column 13   Coefficient 0.03226852
         when "111100011101" => A <= "000000010100110111"; -- Line 242   Column 14   Coefficient 0.00509262
         when "111100011110" => A <= "111111111110110111"; -- Line 242   Column 15   Coefficient -0.00027847
         when "111100011111" => A <= "000000000000000000"; -- Line 242   Column 16   Coefficient 0.00000000
         when "111100100000" => A <= "000000000000000000"; -- Line 243   Column 1   Coefficient 0.00000000
         when "111100100001" => A <= "000000000000000000"; -- Line 243   Column 2   Coefficient 0.00000000
         when "111100100010" => A <= "000000000000000000"; -- Line 243   Column 3   Coefficient 0.00000000
         when "111100100011" => A <= "000000000000000000"; -- Line 243   Column 4   Coefficient 0.00000000
         when "111100100100" => A <= "000000000000000000"; -- Line 243   Column 5   Coefficient 0.00000000
         when "111100100101" => A <= "000000000000000000"; -- Line 243   Column 6   Coefficient 0.00000000
         when "111100100110" => A <= "000000000000000000"; -- Line 243   Column 7   Coefficient 0.00000000
         when "111100100111" => A <= "000000000000000000"; -- Line 243   Column 8   Coefficient 0.00000000
         when "111100101000" => A <= "000000000000000000"; -- Line 243   Column 9   Coefficient 0.00000000
         when "111100101001" => A <= "000000001000010011"; -- Line 243   Column 10   Coefficient 0.00202560
         when "111100101010" => A <= "111101100110110000"; -- Line 243   Column 11   Coefficient -0.03741455
         when "111100101011" => A <= "001110110101010100"; -- Line 243   Column 12   Coefficient 0.23176575
         when "111100101100" => A <= "000011001010010011"; -- Line 243   Column 13   Coefficient 0.04938889
         when "111100101101" => A <= "000000010100111001"; -- Line 243   Column 14   Coefficient 0.00510025
         when "111100101110" => A <= "111111111100011110"; -- Line 243   Column 15   Coefficient -0.00086212
         when "111100101111" => A <= "111111111111111111"; -- Line 243   Column 16   Coefficient -0.00000381
         when "111100110000" => A <= "000000000000000000"; -- Line 244   Column 1   Coefficient 0.00000000
         when "111100110001" => A <= "000000000000000000"; -- Line 244   Column 2   Coefficient 0.00000000
         when "111100110010" => A <= "000000000000000000"; -- Line 244   Column 3   Coefficient 0.00000000
         when "111100110011" => A <= "000000000000000000"; -- Line 244   Column 4   Coefficient 0.00000000
         when "111100110100" => A <= "000000000000000000"; -- Line 244   Column 5   Coefficient 0.00000000
         when "111100110101" => A <= "000000000000000000"; -- Line 244   Column 6   Coefficient 0.00000000
         when "111100110110" => A <= "000000000000000000"; -- Line 244   Column 7   Coefficient 0.00000000
         when "111100110111" => A <= "000000000000000000"; -- Line 244   Column 8   Coefficient 0.00000000
         when "111100111000" => A <= "000000000000000000"; -- Line 244   Column 9   Coefficient 0.00000000
         when "111100111001" => A <= "000000000011111000"; -- Line 244   Column 10   Coefficient 0.00094604
         when "111100111010" => A <= "111101110100001010"; -- Line 244   Column 11   Coefficient -0.03414154
         when "111100111011" => A <= "001101100011111111"; -- Line 244   Column 12   Coefficient 0.21191025
         when "111100111100" => A <= "000100010011001101"; -- Line 244   Column 13   Coefficient 0.06718826
         when "111100111101" => A <= "000000010111101010"; -- Line 244   Column 14   Coefficient 0.00577545
         when "111100111110" => A <= "111111111001000110"; -- Line 244   Column 15   Coefficient -0.00168610
         when "111100111111" => A <= "000000000000000011"; -- Line 244   Column 16   Coefficient 0.00001144
         when "111101000000" => A <= "000000000000000000"; -- Line 245   Column 1   Coefficient 0.00000000
         when "111101000001" => A <= "000000000000000000"; -- Line 245   Column 2   Coefficient 0.00000000
         when "111101000010" => A <= "000000000000000000"; -- Line 245   Column 3   Coefficient 0.00000000
         when "111101000011" => A <= "000000000000000000"; -- Line 245   Column 4   Coefficient 0.00000000
         when "111101000100" => A <= "000000000000000000"; -- Line 245   Column 5   Coefficient 0.00000000
         when "111101000101" => A <= "000000000000000000"; -- Line 245   Column 6   Coefficient 0.00000000
         when "111101000110" => A <= "000000000000000000"; -- Line 245   Column 7   Coefficient 0.00000000
         when "111101000111" => A <= "000000000000000000"; -- Line 245   Column 8   Coefficient 0.00000000
         when "111101001000" => A <= "000000000000000000"; -- Line 245   Column 9   Coefficient 0.00000000
         when "111101001001" => A <= "111111111111010011"; -- Line 245   Column 10   Coefficient -0.00017166
         when "111101001010" => A <= "111110000101010011"; -- Line 245   Column 11   Coefficient -0.02995682
         when "111101001011" => A <= "001100001011101000"; -- Line 245   Column 12   Coefficient 0.19033813
         when "111101001100" => A <= "000101100000010101"; -- Line 245   Column 13   Coefficient 0.08601761
         when "111101001101" => A <= "000000011000110111"; -- Line 245   Column 14   Coefficient 0.00606918
         when "111101001110" => A <= "111111110110011111"; -- Line 245   Column 15   Coefficient -0.00232315
         when "111101001111" => A <= "000000000000000110"; -- Line 245   Column 16   Coefficient 0.00002289
         when "111101010000" => A <= "000000000000000000"; -- Line 246   Column 1   Coefficient 0.00000000
         when "111101010001" => A <= "000000000000000000"; -- Line 246   Column 2   Coefficient 0.00000000
         when "111101010010" => A <= "000000000000000000"; -- Line 246   Column 3   Coefficient 0.00000000
         when "111101010011" => A <= "000000000000000000"; -- Line 246   Column 4   Coefficient 0.00000000
         when "111101010100" => A <= "000000000000000000"; -- Line 246   Column 5   Coefficient 0.00000000
         when "111101010101" => A <= "000000000000000000"; -- Line 246   Column 6   Coefficient 0.00000000
         when "111101010110" => A <= "000000000000000000"; -- Line 246   Column 7   Coefficient 0.00000000
         when "111101010111" => A <= "000000000000000000"; -- Line 246   Column 8   Coefficient 0.00000000
         when "111101011000" => A <= "000000000000000000"; -- Line 246   Column 9   Coefficient 0.00000000
         when "111101011001" => A <= "111111111110010010"; -- Line 246   Column 10   Coefficient -0.00041962
         when "111101011010" => A <= "111110010000110000"; -- Line 246   Column 11   Coefficient -0.02716064
         when "111101011011" => A <= "001010101100000111"; -- Line 246   Column 12   Coefficient 0.16701889
         when "111101011100" => A <= "000111000101010101"; -- Line 246   Column 13   Coefficient 0.11067581
         when "111101011101" => A <= "000000000100100100"; -- Line 246   Column 14   Coefficient 0.00111389
         when "111101011110" => A <= "111111111010111001"; -- Line 246   Column 15   Coefficient -0.00124741
         when "111101011111" => A <= "000000000000000100"; -- Line 246   Column 16   Coefficient 0.00001526
         when "111101100000" => A <= "000000000000000000"; -- Line 247   Column 1   Coefficient 0.00000000
         when "111101100001" => A <= "000000000000000000"; -- Line 247   Column 2   Coefficient 0.00000000
         when "111101100010" => A <= "000000000000000000"; -- Line 247   Column 3   Coefficient 0.00000000
         when "111101100011" => A <= "000000000000000000"; -- Line 247   Column 4   Coefficient 0.00000000
         when "111101100100" => A <= "000000000000000000"; -- Line 247   Column 5   Coefficient 0.00000000
         when "111101100101" => A <= "000000000000000000"; -- Line 247   Column 6   Coefficient 0.00000000
         when "111101100110" => A <= "000000000000000000"; -- Line 247   Column 7   Coefficient 0.00000000
         when "111101100111" => A <= "000000000000000000"; -- Line 247   Column 8   Coefficient 0.00000000
         when "111101101000" => A <= "000000000000000000"; -- Line 247   Column 9   Coefficient 0.00000000
         when "111101101001" => A <= "111111111110100110"; -- Line 247   Column 10   Coefficient -0.00034332
         when "111101101010" => A <= "111110011011111010"; -- Line 247   Column 11   Coefficient -0.02443695
         when "111101101011" => A <= "001001000110101001"; -- Line 247   Column 12   Coefficient 0.14224625
         when "111101101100" => A <= "001000110101000000"; -- Line 247   Column 13   Coefficient 0.13793945
         when "111101101101" => A <= "111111100111100010"; -- Line 247   Column 14   Coefficient -0.00597382
         when "111101101110" => A <= "000000000010010011"; -- Line 247   Column 15   Coefficient 0.00056076
         when "111101101111" => A <= "000000000000000011"; -- Line 247   Column 16   Coefficient 0.00001144
         when "111101110000" => A <= "000000000000000000"; -- Line 248   Column 1   Coefficient 0.00000000
         when "111101110001" => A <= "000000000000000000"; -- Line 248   Column 2   Coefficient 0.00000000
         when "111101110010" => A <= "000000000000000000"; -- Line 248   Column 3   Coefficient 0.00000000
         when "111101110011" => A <= "000000000000000000"; -- Line 248   Column 4   Coefficient 0.00000000
         when "111101110100" => A <= "000000000000000000"; -- Line 248   Column 5   Coefficient 0.00000000
         when "111101110101" => A <= "000000000000000000"; -- Line 248   Column 6   Coefficient 0.00000000
         when "111101110110" => A <= "000000000000000000"; -- Line 248   Column 7   Coefficient 0.00000000
         when "111101110111" => A <= "000000000000000000"; -- Line 248   Column 8   Coefficient 0.00000000
         when "111101111000" => A <= "000000000000000000"; -- Line 248   Column 9   Coefficient 0.00000000
         when "111101111001" => A <= "111111111111001011"; -- Line 248   Column 10   Coefficient -0.00020218
         when "111101111010" => A <= "111110100110010011"; -- Line 248   Column 11   Coefficient -0.02190018
         when "111101111011" => A <= "000111100110110001"; -- Line 248   Column 12   Coefficient 0.11883926
         when "111101111100" => A <= "001010011001111000"; -- Line 248   Column 13   Coefficient 0.16256714
         when "111101111101" => A <= "111111010000101110"; -- Line 248   Column 14   Coefficient -0.01154327
         when "111101111110" => A <= "000000001001011000"; -- Line 248   Column 15   Coefficient 0.00228882
         when "111101111111" => A <= "111111111111110100"; -- Line 248   Column 16   Coefficient -0.00004578
         when "111110000000" => A <= "000000000000000000"; -- Line 249   Column 1   Coefficient 0.00000000
         when "111110000001" => A <= "000000000000000000"; -- Line 249   Column 2   Coefficient 0.00000000
         when "111110000010" => A <= "000000000000000000"; -- Line 249   Column 3   Coefficient 0.00000000
         when "111110000011" => A <= "000000000000000000"; -- Line 249   Column 4   Coefficient 0.00000000
         when "111110000100" => A <= "000000000000000000"; -- Line 249   Column 5   Coefficient 0.00000000
         when "111110000101" => A <= "000000000000000000"; -- Line 249   Column 6   Coefficient 0.00000000
         when "111110000110" => A <= "000000000000000000"; -- Line 249   Column 7   Coefficient 0.00000000
         when "111110000111" => A <= "000000000000000000"; -- Line 249   Column 8   Coefficient 0.00000000
         when "111110001000" => A <= "000000000000000000"; -- Line 249   Column 9   Coefficient 0.00000000
         when "111110001001" => A <= "000000000000000011"; -- Line 249   Column 10   Coefficient 0.00001144
         when "111110001010" => A <= "111110110001100001"; -- Line 249   Column 11   Coefficient -0.01916122
         when "111110001011" => A <= "000110000101110011"; -- Line 249   Column 12   Coefficient 0.09516525
         when "111110001100" => A <= "001011111101111010"; -- Line 249   Column 13   Coefficient 0.18698883
         when "111110001101" => A <= "111110111010000001"; -- Line 249   Column 14   Coefficient -0.01708603
         when "111110001110" => A <= "000000010001001000"; -- Line 249   Column 15   Coefficient 0.00418091
         when "111110001111" => A <= "111111111111100110"; -- Line 249   Column 16   Coefficient -0.00009918
         when "111110010000" => A <= "000000000000000000"; -- Line 250   Column 1   Coefficient 0.00000000
         when "111110010001" => A <= "000000000000000000"; -- Line 250   Column 2   Coefficient 0.00000000
         when "111110010010" => A <= "000000000000000000"; -- Line 250   Column 3   Coefficient 0.00000000
         when "111110010011" => A <= "000000000000000000"; -- Line 250   Column 4   Coefficient 0.00000000
         when "111110010100" => A <= "000000000000000000"; -- Line 250   Column 5   Coefficient 0.00000000
         when "111110010101" => A <= "000000000000000000"; -- Line 250   Column 6   Coefficient 0.00000000
         when "111110010110" => A <= "000000000000000000"; -- Line 250   Column 7   Coefficient 0.00000000
         when "111110010111" => A <= "000000000000000000"; -- Line 250   Column 8   Coefficient 0.00000000
         when "111110011000" => A <= "000000000000000000"; -- Line 250   Column 9   Coefficient 0.00000000
         when "111110011001" => A <= "000000000000001001"; -- Line 250   Column 10   Coefficient 0.00003433
         when "111110011010" => A <= "111111000100111001"; -- Line 250   Column 11   Coefficient -0.01443100
         when "111110011011" => A <= "000100010010000101"; -- Line 250   Column 12   Coefficient 0.06691360
         when "111110011100" => A <= "001101110100101001"; -- Line 250   Column 13   Coefficient 0.21597672
         when "111110011101" => A <= "111110011010010101"; -- Line 250   Column 14   Coefficient -0.02482224
         when "111110011110" => A <= "000000011001110100"; -- Line 250   Column 15   Coefficient 0.00630188
         when "111110011111" => A <= "000000000000000111"; -- Line 250   Column 16   Coefficient 0.00002670
         when "111110100000" => A <= "000000000000000000"; -- Line 251   Column 1   Coefficient 0.00000000
         when "111110100001" => A <= "000000000000000000"; -- Line 251   Column 2   Coefficient 0.00000000
         when "111110100010" => A <= "000000000000000000"; -- Line 251   Column 3   Coefficient 0.00000000
         when "111110100011" => A <= "000000000000000000"; -- Line 251   Column 4   Coefficient 0.00000000
         when "111110100100" => A <= "000000000000000000"; -- Line 251   Column 5   Coefficient 0.00000000
         when "111110100101" => A <= "000000000000000000"; -- Line 251   Column 6   Coefficient 0.00000000
         when "111110100110" => A <= "000000000000000000"; -- Line 251   Column 7   Coefficient 0.00000000
         when "111110100111" => A <= "000000000000000000"; -- Line 251   Column 8   Coefficient 0.00000000
         when "111110101000" => A <= "000000000000000000"; -- Line 251   Column 9   Coefficient 0.00000000
         when "111110101001" => A <= "000000000000000000"; -- Line 251   Column 10   Coefficient 0.00000000
         when "111110101010" => A <= "111111011001111001"; -- Line 251   Column 11   Coefficient -0.00930405
         when "111110101011" => A <= "000010011110111100"; -- Line 251   Column 12   Coefficient 0.03880310
         when "111110101100" => A <= "001111100101110011"; -- Line 251   Column 13   Coefficient 0.24360275
         when "111110101101" => A <= "111101111110110001"; -- Line 251   Column 14   Coefficient -0.03155136
         when "111110101110" => A <= "000000100001110011"; -- Line 251   Column 15   Coefficient 0.00825119
         when "111110101111" => A <= "000000000000110011"; -- Line 251   Column 16   Coefficient 0.00019455
         when "111110110000" => A <= "000000000000000000"; -- Line 252   Column 1   Coefficient 0.00000000
         when "111110110001" => A <= "000000000000000000"; -- Line 252   Column 2   Coefficient 0.00000000
         when "111110110010" => A <= "000000000000000000"; -- Line 252   Column 3   Coefficient 0.00000000
         when "111110110011" => A <= "000000000000000000"; -- Line 252   Column 4   Coefficient 0.00000000
         when "111110110100" => A <= "000000000000000000"; -- Line 252   Column 5   Coefficient 0.00000000
         when "111110110101" => A <= "000000000000000000"; -- Line 252   Column 6   Coefficient 0.00000000
         when "111110110110" => A <= "000000000000000000"; -- Line 252   Column 7   Coefficient 0.00000000
         when "111110110111" => A <= "000000000000000000"; -- Line 252   Column 8   Coefficient 0.00000000
         when "111110111000" => A <= "000000000000000000"; -- Line 252   Column 9   Coefficient 0.00000000
         when "111110111001" => A <= "000000000000000000"; -- Line 252   Column 10   Coefficient 0.00000000
         when "111110111010" => A <= "111111110001010101"; -- Line 252   Column 11   Coefficient -0.00358200
         when "111110111011" => A <= "000000100101011001"; -- Line 252   Column 12   Coefficient 0.00912857
         when "111110111100" => A <= "010001011110001011"; -- Line 252   Column 13   Coefficient 0.27299118
         when "111110111101" => A <= "111101011101101101"; -- Line 252   Column 14   Coefficient -0.03962326
         when "111110111110" => A <= "000000101011110101"; -- Line 252   Column 15   Coefficient 0.01070023
         when "111110111111" => A <= "000000000001100101"; -- Line 252   Column 16   Coefficient 0.00038528
         when "111111000000" => A <= "000000000000000000"; -- Line 253   Column 1   Coefficient 0.00000000
         when "111111000001" => A <= "000000000000000000"; -- Line 253   Column 2   Coefficient 0.00000000
         when "111111000010" => A <= "000000000000000000"; -- Line 253   Column 3   Coefficient 0.00000000
         when "111111000011" => A <= "000000000000000000"; -- Line 253   Column 4   Coefficient 0.00000000
         when "111111000100" => A <= "000000000000000000"; -- Line 253   Column 5   Coefficient 0.00000000
         when "111111000101" => A <= "000000000000000000"; -- Line 253   Column 6   Coefficient 0.00000000
         when "111111000110" => A <= "000000000000000000"; -- Line 253   Column 7   Coefficient 0.00000000
         when "111111000111" => A <= "000000000000000000"; -- Line 253   Column 8   Coefficient 0.00000000
         when "111111001000" => A <= "000000000000000000"; -- Line 253   Column 9   Coefficient 0.00000000
         when "111111001001" => A <= "000000000000000000"; -- Line 253   Column 10   Coefficient 0.00000000
         when "111111001010" => A <= "000000000111011010"; -- Line 253   Column 11   Coefficient 0.00180817
         when "111111001011" => A <= "111110110101100100"; -- Line 253   Column 12   Coefficient -0.01817322
         when "111111001100" => A <= "010011000101100111"; -- Line 253   Column 13   Coefficient 0.29824448
         when "111111001101" => A <= "111101000110110001"; -- Line 253   Column 14   Coefficient -0.04522324
         when "111111001110" => A <= "000000110100010110"; -- Line 253   Column 15   Coefficient 0.01277924
         when "111111001111" => A <= "000000000010010101"; -- Line 253   Column 16   Coefficient 0.00056839
         when "111111010000" => A <= "000000000000000000"; -- Line 254   Column 1   Coefficient 0.00000000
         when "111111010001" => A <= "000000000000000000"; -- Line 254   Column 2   Coefficient 0.00000000
         when "111111010010" => A <= "000000000000000000"; -- Line 254   Column 3   Coefficient 0.00000000
         when "111111010011" => A <= "000000000000000000"; -- Line 254   Column 4   Coefficient 0.00000000
         when "111111010100" => A <= "000000000000000000"; -- Line 254   Column 5   Coefficient 0.00000000
         when "111111010101" => A <= "000000000000000000"; -- Line 254   Column 6   Coefficient 0.00000000
         when "111111010110" => A <= "000000000000000000"; -- Line 254   Column 7   Coefficient 0.00000000
         when "111111010111" => A <= "000000000000000000"; -- Line 254   Column 8   Coefficient 0.00000000
         when "111111011000" => A <= "000000000000000000"; -- Line 254   Column 9   Coefficient 0.00000000
         when "111111011001" => A <= "000000000000000000"; -- Line 254   Column 10   Coefficient 0.00000000
         when "111111011010" => A <= "000000001111000010"; -- Line 254   Column 11   Coefficient 0.00366974
         when "111111011011" => A <= "111110000010011110"; -- Line 254   Column 12   Coefficient -0.03064728
         when "111111011100" => A <= "010011010010100110"; -- Line 254   Column 13   Coefficient 0.30141449
         when "111111011101" => A <= "111101100111001110"; -- Line 254   Column 14   Coefficient -0.03730011
         when "111111011110" => A <= "000000110010101110"; -- Line 254   Column 15   Coefficient 0.01238251
         when "111111011111" => A <= "000000000001111110"; -- Line 254   Column 16   Coefficient 0.00048065
         when "111111100000" => A <= "000000000000000000"; -- Line 255   Column 1   Coefficient 0.00000000
         when "111111100001" => A <= "000000000000000000"; -- Line 255   Column 2   Coefficient 0.00000000
         when "111111100010" => A <= "000000000000000000"; -- Line 255   Column 3   Coefficient 0.00000000
         when "111111100011" => A <= "000000000000000000"; -- Line 255   Column 4   Coefficient 0.00000000
         when "111111100100" => A <= "000000000000000000"; -- Line 255   Column 5   Coefficient 0.00000000
         when "111111100101" => A <= "000000000000000000"; -- Line 255   Column 6   Coefficient 0.00000000
         when "111111100110" => A <= "000000000000000000"; -- Line 255   Column 7   Coefficient 0.00000000
         when "111111100111" => A <= "000000000000000000"; -- Line 255   Column 8   Coefficient 0.00000000
         when "111111101000" => A <= "000000000000000000"; -- Line 255   Column 9   Coefficient 0.00000000
         when "111111101001" => A <= "000000000000000000"; -- Line 255   Column 10   Coefficient 0.00000000
         when "111111101010" => A <= "000000010000011000"; -- Line 255   Column 11   Coefficient 0.00399780
         when "111111101011" => A <= "111101101011101110"; -- Line 255   Column 12   Coefficient -0.03620148
         when "111111101100" => A <= "010010110100110100"; -- Line 255   Column 13   Coefficient 0.29414368
         when "111111101101" => A <= "111110100000101100"; -- Line 255   Column 14   Coefficient -0.02326965
         when "111111101110" => A <= "000000101101010111"; -- Line 255   Column 15   Coefficient 0.01107407
         when "111111101111" => A <= "000000000001000010"; -- Line 255   Column 16   Coefficient 0.00025177
         when "111111110000" => A <= "000000000000000000"; -- Line 256   Column 1   Coefficient 0.00000000
         when "111111110001" => A <= "000000000000000000"; -- Line 256   Column 2   Coefficient 0.00000000
         when "111111110010" => A <= "000000000000000000"; -- Line 256   Column 3   Coefficient 0.00000000
         when "111111110011" => A <= "000000000000000000"; -- Line 256   Column 4   Coefficient 0.00000000
         when "111111110100" => A <= "000000000000000000"; -- Line 256   Column 5   Coefficient 0.00000000
         when "111111110101" => A <= "000000000000000000"; -- Line 256   Column 6   Coefficient 0.00000000
         when "111111110110" => A <= "000000000000000000"; -- Line 256   Column 7   Coefficient 0.00000000
         when "111111110111" => A <= "000000000000000000"; -- Line 256   Column 8   Coefficient 0.00000000
         when "111111111000" => A <= "000000000000000000"; -- Line 256   Column 9   Coefficient 0.00000000
         when "111111111001" => A <= "000000000000000000"; -- Line 256   Column 10   Coefficient 0.00000000
         when "111111111010" => A <= "000000001111111100"; -- Line 256   Column 11   Coefficient 0.00389099
         when "111111111011" => A <= "111101100000101101"; -- Line 256   Column 12   Coefficient -0.03889084
         when "111111111100" => A <= "010010000001100011"; -- Line 256   Column 13   Coefficient 0.28162766
         when "111111111101" => A <= "111111101010001000"; -- Line 256   Column 14   Coefficient -0.00534058
         when "111111111110" => A <= "000000100010100100"; -- Line 256   Column 15   Coefficient 0.00843811
         when "111111111111" => A <= "000000000001001000"; -- Line 256   Column 16   Coefficient 0.00027466
         when others => null;
      end case;
   end process;
end LUTable;
