library ieee;
use ieee.std_logic_1164.all;

entity fsm_toggle is

	generic(
	
	n :	integer := 4
	
	);

	port(
	
	RST,CLK : in std_logic;
	
	pmt : in std_logic;
	
	bt_sample : in std_logic;
	bt_window : in std_logic;
	bt_int : in std_logic;
	bt_n : in std_logic;
	
	clr_sample : out std_logic;
	clr_window : out std_logic;
	clr_int : out std_logic;
	clr_n : out std_logic;
	
	adc_clk : out std_logic;
	int_rst : out std_logic;
	data_valid : out std_logic;
	sample_c : out std_logic
	
	);
end fsm_toggle;

architecture fsm of fsm_toggle is	


signal qp, qn : std_logic_vector(n-1 downto 0);

begin  
	
	c1 : process(qp,pmt,bt_sample,bt_int,bt_window,bt_n)
	begin
		
		case(qp) is
		
		--s0
		when "0000" =>
		clr_sample <= '1'; 
		clr_window <= '1';
		clr_int <= '1';
		clr_n <= '1';
		adc_clk <= '0';
		int_rst <= '1';
		data_valid <= '0';
		sample_c <= '0';
		
		if(pmt='1') then
			qn <= "0001";
		else
			qn <= "0000";
		end if;
		
		--s1
		when "0001" =>
		clr_sample <= '0';
		clr_window <= '0';	
		clr_int <= '0';
		clr_n <= '1';
		adc_clk <= '0';
		int_rst <= '0';   --ventana de integracion
		data_valid <= '0';
		sample_c <= '0';
		
		if(bt_int='1') then
			qn <= "0010";
		else
			qn <= "0001";
		end if;
		
		--s2
		when "0010" =>
		clr_sample <= '0';
		clr_window <= '0';	
		clr_int <= '0';
		clr_n <= '1';
		adc_clk <= '1';
		int_rst <= '0';   --ventana de integracion
		data_valid <= '0';
		sample_c <= '0';
		
		if(bt_window='1') then
			qn <= "0011";
		else
			qn <= "0010";
		end if;
		
		--s3 subes 1
		when "0011" =>
		clr_sample <= '0';
		clr_window <= '0';	
		clr_int <= '1';
		clr_n <= '0';
		adc_clk <= '1';
		int_rst <= '1';   --reset integragor
		data_valid <= '0';
		sample_c <= '0';
		
		if(bt_n='1') then
			qn <= "0100";
		else
			qn <= "0011";
		end if;
		
		--s4 bajas
		when "0100" =>
		clr_sample <= '0';
		clr_window <= '1';	
		clr_int <= '1';
		clr_n <= '0';
		adc_clk <= '0';
		int_rst <= '1';   --reset integragor
		data_valid <= '0';
		sample_c <= '0';
		
		if(bt_n='1') then
			qn <= "0101";
		else
			qn <= "0100";
		end if;
		
		--s5 subes 2
		when "0101" =>
		clr_sample <= '0';
		clr_window <= '1';	
		clr_int <= '1';
		clr_n <= '0';
		adc_clk <= '1';
		int_rst <= '1';   --reset integragor
		data_valid <= '0';
		sample_c <= '0';
		
		if(bt_n='1') then
			qn <= "0110";
		else
			qn <= "0101";
		end if;
		
		--s6 bajas
		when "0110" =>
		clr_sample <= '0';
		clr_window <= '1';	
		clr_int <= '1';
		clr_n <= '0';
		adc_clk <= '0';
		int_rst <= '1';   --reset integragor
		data_valid <= '0';
		sample_c <= '0';
		
		if(bt_n='1') then
			qn <= "0111";
		else
			qn <= "0110";
		end if;
		
		--s7 subes 3
		when "0111" =>
		clr_sample <= '0';
		clr_window <= '1';	
		clr_int <= '1';
		clr_n <= '0';
		adc_clk <= '1';
		int_rst <= '1';   --reset integragor
		data_valid <= '0';
		sample_c <= '0';
		
		if(bt_n='1') then
			qn <= "1000";
		else
			qn <= "0111";
		end if;
		
		--s8 bajas 
		when "1000" =>
		clr_sample <= '0';
		clr_window <= '1';	
		clr_int <= '1';
		clr_n <= '0';
		adc_clk <= '0';
		int_rst <= '1';   --reset integragor
		data_valid <= '0';
		sample_c <= '0';
		
		if(bt_n='1') then
			qn <= "1001";
		else
			qn <= "1000";
		end if;
		
		
		--s9 subes 4
		when "1001" =>
		clr_sample <= '0';
		clr_window <= '1';	
		clr_int <= '1';
		clr_n <= '0';
		adc_clk <= '1';
		int_rst <= '1';   --reset integragor
		data_valid <= '0';
		sample_c <= '0';
		
		if(bt_n='1') then
			qn <= "1010";
		else
			qn <= "1001";
		end if;
		
		--s10 bajas
		when "1010" =>
		clr_sample <= '0';
		clr_window <= '1';	
		clr_int <= '1';
		clr_n <= '0';
		adc_clk <= '0';
		int_rst <= '1';   --reset integragor
		data_valid <= '0';
		sample_c <= '0';
		
		if(bt_n='1') then
			qn <= "1011";
		else
			qn <= "1010";
		end if;
		
		--s11
		when "1011" =>
		clr_sample <= '0';
		clr_window <= '1';	
		clr_int <= '1';
		clr_n <= '0';
		adc_clk <= '0';
		int_rst <= '1';   --reset integragor
		data_valid <= '0';
		sample_c <= '0';
		
		if(bt_n='1') then
			qn <= "1100";
		else
			qn <= "1011";
		end if;
		
		--s12
		when "1100" =>
		clr_sample <= '0';
		clr_window <= '1';	
		clr_int <= '1';
		clr_n <= '1';
		adc_clk <= '0';
		int_rst <= '1';   --reset integragor
		data_valid <= '1';  --valid
		sample_c <= '0';
		
		qn <= "1101";
		
		--s13
		when "1101" =>
		clr_sample <= '0';
		clr_window <= '1';	
		clr_int <= '1';
		clr_n <= '1';
		adc_clk <= '0';
		int_rst <= '1';   --reset integragor
		data_valid <= '0';
		sample_c <= '0';
		
		qn <= "1110";
		
		--s14
		when "1110" =>
		clr_sample <= '0';
		clr_window <= '1';	
		clr_int <= '1';
		clr_n <= '1';
		adc_clk <= '0';
		int_rst <= '1';   --reset integragor
		data_valid <= '0'; 
		sample_c <= '1';  --counter sample
		
		qn <= "1111";
		
		--s15
		when others =>
		clr_sample <= '0';
		clr_window <= '1';	
		clr_int <= '1';
		clr_n <= '1';
		adc_clk <= '0';
		int_rst <= '1';   --reset integragor
		data_valid <= '0'; 
		sample_c <= '0'; 
		
		if(bt_sample='1') then
			qn <= "0000";
		else
			qn <= "1111";
		end if;
	
		end case;
		
	end process;
	
	secuencial : process(RST,CLK)
	begin
		if(RST='0') then
			qp <= (others => '0');
		elsif(CLK'event and CLK='1') then
			qp <= qn;
		end if;
	end process;
	
end fsm;