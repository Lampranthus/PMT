library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM_20LOG10 is
   port(
      CLK : in std_logic;
      I   : in  std_logic_vector(11 downto 0);
      A   : out std_logic_vector(17 downto 0)
      );
   end ROM_20LOG10;

architecture ROM of ROM_20LOG10 is

subtype word_t is std_logic_vector(17 downto 0);
type memory_t is array(0 to 4095) of word_t;

signal rom : memory_t := (         -- Coefficient format 8.10
   "000000000000000000", -- Line 1   Column 1   Coefficient 0.00000000
   "000001100000010101", -- Line 1   Column 2   Coefficient 6.02050781
   "000010011000101011", -- Line 1   Column 3   Coefficient 9.54199219
   "000011000000101010", -- Line 1   Column 4   Coefficient 12.04101563
   "000011011111101011", -- Line 1   Column 5   Coefficient 13.97949219
   "000011111001000001", -- Line 1   Column 6   Coefficient 15.56347656
   "000100001110011100", -- Line 1   Column 7   Coefficient 16.90234375
   "000100100000111111", -- Line 1   Column 8   Coefficient 18.06152344
   "000100110001010111", -- Line 1   Column 9   Coefficient 19.08496094
   "000101000000000000", -- Line 1   Column 10   Coefficient 20.00000000
   "000101001101010000", -- Line 1   Column 11   Coefficient 20.82812500
   "000101011001010110", -- Line 1   Column 12   Coefficient 21.58398438
   "000101100100011110", -- Line 1   Column 13   Coefficient 22.27929688
   "000101101110110001", -- Line 1   Column 14   Coefficient 22.92285156
   "000101111000010110", -- Line 1   Column 15   Coefficient 23.52148438
   "000110000001010100", -- Line 1   Column 16   Coefficient 24.08203125
   "000110001001110000", -- Line 1   Column 17   Coefficient 24.60937500
   "000110010001101100", -- Line 1   Column 18   Coefficient 25.10546875
   "000110011001001101", -- Line 1   Column 19   Coefficient 25.57519531
   "000110100000010101", -- Line 1   Column 20   Coefficient 26.02050781
   "000110100111000111", -- Line 1   Column 21   Coefficient 26.44433594
   "000110101101100101", -- Line 1   Column 22   Coefficient 26.84863281
   "000110110011110000", -- Line 1   Column 23   Coefficient 27.23437500
   "000110111001101011", -- Line 1   Column 24   Coefficient 27.60449219
   "000110111111010110", -- Line 1   Column 25   Coefficient 27.95898438
   "000111000100110011", -- Line 1   Column 26   Coefficient 28.29980469
   "000111001010000010", -- Line 1   Column 27   Coefficient 28.62695313
   "000111001111000110", -- Line 1   Column 28   Coefficient 28.94335938
   "000111010011111110", -- Line 1   Column 29   Coefficient 29.24804688
   "000111011000101011", -- Line 1   Column 30   Coefficient 29.54199219
   "000111011101001111", -- Line 1   Column 31   Coefficient 29.82714844
   "000111100001101001", -- Line 1   Column 32   Coefficient 30.10253906
   "000111100101111011", -- Line 1   Column 33   Coefficient 30.37011719
   "000111101010000101", -- Line 1   Column 34   Coefficient 30.62988281
   "000111101110000111", -- Line 1   Column 35   Coefficient 30.88183594
   "000111110010000001", -- Line 1   Column 36   Coefficient 31.12597656
   "000111110101110101", -- Line 1   Column 37   Coefficient 31.36425781
   "000111111001100010", -- Line 1   Column 38   Coefficient 31.59570313
   "000111111101001001", -- Line 1   Column 39   Coefficient 31.82128906
   "001000000000101010", -- Line 1   Column 40   Coefficient 32.04101563
   "001000000100000110", -- Line 1   Column 41   Coefficient 32.25585938
   "001000000111011100", -- Line 1   Column 42   Coefficient 32.46484375
   "001000001010101101", -- Line 1   Column 43   Coefficient 32.66894531
   "001000001101111010", -- Line 1   Column 44   Coefficient 32.86914063
   "001000010001000010", -- Line 1   Column 45   Coefficient 33.06445313
   "001000010100000101", -- Line 1   Column 46   Coefficient 33.25488281
   "001000010111000101", -- Line 1   Column 47   Coefficient 33.44238281
   "001000011010000000", -- Line 1   Column 48   Coefficient 33.62500000
   "001000011100110111", -- Line 1   Column 49   Coefficient 33.80371094
   "001000011111101011", -- Line 1   Column 50   Coefficient 33.97949219
   "001000100010011011", -- Line 1   Column 51   Coefficient 34.15136719
   "001000100101001000", -- Line 1   Column 52   Coefficient 34.32031250
   "001000100111110001", -- Line 1   Column 53   Coefficient 34.48535156
   "001000101010010111", -- Line 1   Column 54   Coefficient 34.64746094
   "001000101100111011", -- Line 1   Column 55   Coefficient 34.80761719
   "001000101111011011", -- Line 1   Column 56   Coefficient 34.96386719
   "001000110001111000", -- Line 1   Column 57   Coefficient 35.11718750
   "001000110100010011", -- Line 1   Column 58   Coefficient 35.26855469
   "001000110110101011", -- Line 1   Column 59   Coefficient 35.41699219
   "001000111001000001", -- Line 1   Column 60   Coefficient 35.56347656
   "001000111011010100", -- Line 1   Column 61   Coefficient 35.70703125
   "001000111101100100", -- Line 1   Column 62   Coefficient 35.84765625
   "001000111111110010", -- Line 1   Column 63   Coefficient 35.98632813
   "001001000001111111", -- Line 1   Column 64   Coefficient 36.12402344
   "001001000100001000", -- Line 1   Column 65   Coefficient 36.25781250
   "001001000110010000", -- Line 1   Column 66   Coefficient 36.39062500
   "001001001000010110", -- Line 1   Column 67   Coefficient 36.52148438
   "001001001010011010", -- Line 1   Column 68   Coefficient 36.65039063
   "001001001100011100", -- Line 1   Column 69   Coefficient 36.77734375
   "001001001110011100", -- Line 1   Column 70   Coefficient 36.90234375
   "001001010000011010", -- Line 1   Column 71   Coefficient 37.02539063
   "001001010010010110", -- Line 1   Column 72   Coefficient 37.14648438
   "001001010100010001", -- Line 1   Column 73   Coefficient 37.26660156
   "001001010110001010", -- Line 1   Column 74   Coefficient 37.38476563
   "001001011000000001", -- Line 1   Column 75   Coefficient 37.50097656
   "001001011001110111", -- Line 1   Column 76   Coefficient 37.61621094
   "001001011011101011", -- Line 1   Column 77   Coefficient 37.72949219
   "001001011101011110", -- Line 1   Column 78   Coefficient 37.84179688
   "001001011111001111", -- Line 1   Column 79   Coefficient 37.95214844
   "001001100000111111", -- Line 1   Column 80   Coefficient 38.06152344
   "001001100010101110", -- Line 1   Column 81   Coefficient 38.16992188
   "001001100100011011", -- Line 1   Column 82   Coefficient 38.27636719
   "001001100110000111", -- Line 1   Column 83   Coefficient 38.38183594
   "001001100111110001", -- Line 1   Column 84   Coefficient 38.48535156
   "001001101001011010", -- Line 1   Column 85   Coefficient 38.58789063
   "001001101011000011", -- Line 1   Column 86   Coefficient 38.69042969
   "001001101100101001", -- Line 1   Column 87   Coefficient 38.79003906
   "001001101110001111", -- Line 1   Column 88   Coefficient 38.88964844
   "001001101111110100", -- Line 1   Column 89   Coefficient 38.98828125
   "001001110001010111", -- Line 1   Column 90   Coefficient 39.08496094
   "001001110010111001", -- Line 1   Column 91   Coefficient 39.18066406
   "001001110100011010", -- Line 1   Column 92   Coefficient 39.27539063
   "001001110101111011", -- Line 1   Column 93   Coefficient 39.37011719
   "001001110111011010", -- Line 1   Column 94   Coefficient 39.46289063
   "001001111000111000", -- Line 1   Column 95   Coefficient 39.55468750
   "001001111010010101", -- Line 1   Column 96   Coefficient 39.64550781
   "001001111011110001", -- Line 1   Column 97   Coefficient 39.73535156
   "001001111101001100", -- Line 1   Column 98   Coefficient 39.82421875
   "001001111110100111", -- Line 1   Column 99   Coefficient 39.91308594
   "001010000000000000", -- Line 1   Column 100   Coefficient 40.00000000
   "001010000001011001", -- Line 1   Column 101   Coefficient 40.08691406
   "001010000010110000", -- Line 1   Column 102   Coefficient 40.17187500
   "001010000100000111", -- Line 1   Column 103   Coefficient 40.25683594
   "001010000101011101", -- Line 1   Column 104   Coefficient 40.34082031
   "001010000110110010", -- Line 1   Column 105   Coefficient 40.42382813
   "001010001000000110", -- Line 1   Column 106   Coefficient 40.50585938
   "001010001001011010", -- Line 1   Column 107   Coefficient 40.58789063
   "001010001010101101", -- Line 1   Column 108   Coefficient 40.66894531
   "001010001011111110", -- Line 1   Column 109   Coefficient 40.74804688
   "001010001101010000", -- Line 1   Column 110   Coefficient 40.82812500
   "001010001110100000", -- Line 1   Column 111   Coefficient 40.90625000
   "001010001111110000", -- Line 1   Column 112   Coefficient 40.98437500
   "001010010000111111", -- Line 1   Column 113   Coefficient 41.06152344
   "001010010010001101", -- Line 1   Column 114   Coefficient 41.13769531
   "001010010011011011", -- Line 1   Column 115   Coefficient 41.21386719
   "001010010100101000", -- Line 1   Column 116   Coefficient 41.28906250
   "001010010101110100", -- Line 1   Column 117   Coefficient 41.36328125
   "001010010111000000", -- Line 1   Column 118   Coefficient 41.43750000
   "001010011000001011", -- Line 1   Column 119   Coefficient 41.51074219
   "001010011001010110", -- Line 1   Column 120   Coefficient 41.58398438
   "001010011010011111", -- Line 1   Column 121   Coefficient 41.65527344
   "001010011011101001", -- Line 1   Column 122   Coefficient 41.72753906
   "001010011100110001", -- Line 1   Column 123   Coefficient 41.79785156
   "001010011101111001", -- Line 1   Column 124   Coefficient 41.86816406
   "001010011111000001", -- Line 1   Column 125   Coefficient 41.93847656
   "001010100000001000", -- Line 1   Column 126   Coefficient 42.00781250
   "001010100001001110", -- Line 1   Column 127   Coefficient 42.07617188
   "001010100010010100", -- Line 1   Column 128   Coefficient 42.14453125
   "001010100011011001", -- Line 1   Column 129   Coefficient 42.21191406
   "001010100100011110", -- Line 1   Column 130   Coefficient 42.27929688
   "001010100101100010", -- Line 1   Column 131   Coefficient 42.34570313
   "001010100110100101", -- Line 1   Column 132   Coefficient 42.41113281
   "001010100111101000", -- Line 1   Column 133   Coefficient 42.47656250
   "001010101000101011", -- Line 1   Column 134   Coefficient 42.54199219
   "001010101001101101", -- Line 1   Column 135   Coefficient 42.60644531
   "001010101010101111", -- Line 1   Column 136   Coefficient 42.67089844
   "001010101011110000", -- Line 1   Column 137   Coefficient 42.73437500
   "001010101100110001", -- Line 1   Column 138   Coefficient 42.79785156
   "001010101101110001", -- Line 1   Column 139   Coefficient 42.86035156
   "001010101110110001", -- Line 1   Column 140   Coefficient 42.92285156
   "001010101111110000", -- Line 1   Column 141   Coefficient 42.98437500
   "001010110000101111", -- Line 1   Column 142   Coefficient 43.04589844
   "001010110001101101", -- Line 1   Column 143   Coefficient 43.10644531
   "001010110010101011", -- Line 1   Column 144   Coefficient 43.16699219
   "001010110011101001", -- Line 1   Column 145   Coefficient 43.22753906
   "001010110100100110", -- Line 1   Column 146   Coefficient 43.28710938
   "001010110101100011", -- Line 1   Column 147   Coefficient 43.34667969
   "001010110110011111", -- Line 1   Column 148   Coefficient 43.40527344
   "001010110111011011", -- Line 1   Column 149   Coefficient 43.46386719
   "001010111000010110", -- Line 1   Column 150   Coefficient 43.52148438
   "001010111001010001", -- Line 1   Column 151   Coefficient 43.57910156
   "001010111010001100", -- Line 1   Column 152   Coefficient 43.63671875
   "001010111011000110", -- Line 1   Column 153   Coefficient 43.69335938
   "001010111100000000", -- Line 1   Column 154   Coefficient 43.75000000
   "001010111100111010", -- Line 1   Column 155   Coefficient 43.80664063
   "001010111101110011", -- Line 1   Column 156   Coefficient 43.86230469
   "001010111110101100", -- Line 1   Column 157   Coefficient 43.91796875
   "001010111111100100", -- Line 1   Column 158   Coefficient 43.97265625
   "001011000000011101", -- Line 1   Column 159   Coefficient 44.02832031
   "001011000001010100", -- Line 1   Column 160   Coefficient 44.08203125
   "001011000010001100", -- Line 1   Column 161   Coefficient 44.13671875
   "001011000011000011", -- Line 1   Column 162   Coefficient 44.19042969
   "001011000011111010", -- Line 1   Column 163   Coefficient 44.24414063
   "001011000100110000", -- Line 1   Column 164   Coefficient 44.29687500
   "001011000101100110", -- Line 1   Column 165   Coefficient 44.34960938
   "001011000110011100", -- Line 1   Column 166   Coefficient 44.40234375
   "001011000111010001", -- Line 1   Column 167   Coefficient 44.45410156
   "001011001000000110", -- Line 1   Column 168   Coefficient 44.50585938
   "001011001000111011", -- Line 1   Column 169   Coefficient 44.55761719
   "001011001001110000", -- Line 1   Column 170   Coefficient 44.60937500
   "001011001010100100", -- Line 1   Column 171   Coefficient 44.66015625
   "001011001011011000", -- Line 1   Column 172   Coefficient 44.71093750
   "001011001100001011", -- Line 1   Column 173   Coefficient 44.76074219
   "001011001100111110", -- Line 1   Column 174   Coefficient 44.81054688
   "001011001101110001", -- Line 1   Column 175   Coefficient 44.86035156
   "001011001110100100", -- Line 1   Column 176   Coefficient 44.91015625
   "001011001111010110", -- Line 1   Column 177   Coefficient 44.95898438
   "001011010000001001", -- Line 1   Column 178   Coefficient 45.00878906
   "001011010000111010", -- Line 1   Column 179   Coefficient 45.05664063
   "001011010001101100", -- Line 1   Column 180   Coefficient 45.10546875
   "001011010010011101", -- Line 1   Column 181   Coefficient 45.15332031
   "001011010011001110", -- Line 1   Column 182   Coefficient 45.20117188
   "001011010011111111", -- Line 1   Column 183   Coefficient 45.24902344
   "001011010100101111", -- Line 1   Column 184   Coefficient 45.29589844
   "001011010101100000", -- Line 1   Column 185   Coefficient 45.34375000
   "001011010110010000", -- Line 1   Column 186   Coefficient 45.39062500
   "001011010110111111", -- Line 1   Column 187   Coefficient 45.43652344
   "001011010111101111", -- Line 1   Column 188   Coefficient 45.48339844
   "001011011000011110", -- Line 1   Column 189   Coefficient 45.52929688
   "001011011001001101", -- Line 1   Column 190   Coefficient 45.57519531
   "001011011001111100", -- Line 1   Column 191   Coefficient 45.62109375
   "001011011010101010", -- Line 1   Column 192   Coefficient 45.66601563
   "001011011011011000", -- Line 1   Column 193   Coefficient 45.71093750
   "001011011100000110", -- Line 1   Column 194   Coefficient 45.75585938
   "001011011100110100", -- Line 1   Column 195   Coefficient 45.80078125
   "001011011101100001", -- Line 1   Column 196   Coefficient 45.84472656
   "001011011110001111", -- Line 1   Column 197   Coefficient 45.88964844
   "001011011110111100", -- Line 1   Column 198   Coefficient 45.93359375
   "001011011111101001", -- Line 1   Column 199   Coefficient 45.97753906
   "001011100000010101", -- Line 1   Column 200   Coefficient 46.02050781
   "001011100001000001", -- Line 1   Column 201   Coefficient 46.06347656
   "001011100001101110", -- Line 1   Column 202   Coefficient 46.10742188
   "001011100010011010", -- Line 1   Column 203   Coefficient 46.15039063
   "001011100011000101", -- Line 1   Column 204   Coefficient 46.19238281
   "001011100011110001", -- Line 1   Column 205   Coefficient 46.23535156
   "001011100100011100", -- Line 1   Column 206   Coefficient 46.27734375
   "001011100101000111", -- Line 1   Column 207   Coefficient 46.31933594
   "001011100101110010", -- Line 1   Column 208   Coefficient 46.36132813
   "001011100110011101", -- Line 1   Column 209   Coefficient 46.40332031
   "001011100111000111", -- Line 1   Column 210   Coefficient 46.44433594
   "001011100111110001", -- Line 1   Column 211   Coefficient 46.48535156
   "001011101000011011", -- Line 1   Column 212   Coefficient 46.52636719
   "001011101001000101", -- Line 1   Column 213   Coefficient 46.56738281
   "001011101001101111", -- Line 1   Column 214   Coefficient 46.60839844
   "001011101010011000", -- Line 1   Column 215   Coefficient 46.64843750
   "001011101011000010", -- Line 1   Column 216   Coefficient 46.68945313
   "001011101011101011", -- Line 1   Column 217   Coefficient 46.72949219
   "001011101100010100", -- Line 1   Column 218   Coefficient 46.76953125
   "001011101100111100", -- Line 1   Column 219   Coefficient 46.80859375
   "001011101101100101", -- Line 1   Column 220   Coefficient 46.84863281
   "001011101110001101", -- Line 1   Column 221   Coefficient 46.88769531
   "001011101110110101", -- Line 1   Column 222   Coefficient 46.92675781
   "001011101111011101", -- Line 1   Column 223   Coefficient 46.96582031
   "001011110000000101", -- Line 1   Column 224   Coefficient 47.00488281
   "001011110000101101", -- Line 1   Column 225   Coefficient 47.04394531
   "001011110001010100", -- Line 1   Column 226   Coefficient 47.08203125
   "001011110001111011", -- Line 1   Column 227   Coefficient 47.12011719
   "001011110010100011", -- Line 1   Column 228   Coefficient 47.15917969
   "001011110011001001", -- Line 1   Column 229   Coefficient 47.19628906
   "001011110011110000", -- Line 1   Column 230   Coefficient 47.23437500
   "001011110100010111", -- Line 1   Column 231   Coefficient 47.27246094
   "001011110100111101", -- Line 1   Column 232   Coefficient 47.30957031
   "001011110101100011", -- Line 1   Column 233   Coefficient 47.34667969
   "001011110110001010", -- Line 1   Column 234   Coefficient 47.38476563
   "001011110110101111", -- Line 1   Column 235   Coefficient 47.42089844
   "001011110111010101", -- Line 1   Column 236   Coefficient 47.45800781
   "001011110111111011", -- Line 1   Column 237   Coefficient 47.49511719
   "001011111000100000", -- Line 1   Column 238   Coefficient 47.53125000
   "001011111001000110", -- Line 1   Column 239   Coefficient 47.56835938
   "001011111001101011", -- Line 1   Column 240   Coefficient 47.60449219
   "001011111010010000", -- Line 1   Column 241   Coefficient 47.64062500
   "001011111010110101", -- Line 1   Column 242   Coefficient 47.67675781
   "001011111011011001", -- Line 1   Column 243   Coefficient 47.71191406
   "001011111011111110", -- Line 1   Column 244   Coefficient 47.74804688
   "001011111100100010", -- Line 1   Column 245   Coefficient 47.78320313
   "001011111101000110", -- Line 1   Column 246   Coefficient 47.81835938
   "001011111101101010", -- Line 1   Column 247   Coefficient 47.85351563
   "001011111110001110", -- Line 1   Column 248   Coefficient 47.88867188
   "001011111110110010", -- Line 1   Column 249   Coefficient 47.92382813
   "001011111111010110", -- Line 1   Column 250   Coefficient 47.95898438
   "001011111111111001", -- Line 1   Column 251   Coefficient 47.99316406
   "001100000000011101", -- Line 1   Column 252   Coefficient 48.02832031
   "001100000001000000", -- Line 1   Column 253   Coefficient 48.06250000
   "001100000001100011", -- Line 1   Column 254   Coefficient 48.09667969
   "001100000010000110", -- Line 1   Column 255   Coefficient 48.13085938
   "001100000010101001", -- Line 1   Column 256   Coefficient 48.16503906
   "001100000011001011", -- Line 1   Column 257   Coefficient 48.19824219
   "001100000011101110", -- Line 1   Column 258   Coefficient 48.23242188
   "001100000100010000", -- Line 1   Column 259   Coefficient 48.26562500
   "001100000100110011", -- Line 1   Column 260   Coefficient 48.29980469
   "001100000101010101", -- Line 1   Column 261   Coefficient 48.33300781
   "001100000101110111", -- Line 1   Column 262   Coefficient 48.36621094
   "001100000110011001", -- Line 1   Column 263   Coefficient 48.39941406
   "001100000110111010", -- Line 1   Column 264   Coefficient 48.43164063
   "001100000111011100", -- Line 1   Column 265   Coefficient 48.46484375
   "001100000111111110", -- Line 1   Column 266   Coefficient 48.49804688
   "001100001000011111", -- Line 1   Column 267   Coefficient 48.53027344
   "001100001001000000", -- Line 1   Column 268   Coefficient 48.56250000
   "001100001001100001", -- Line 1   Column 269   Coefficient 48.59472656
   "001100001010000010", -- Line 1   Column 270   Coefficient 48.62695313
   "001100001010100011", -- Line 1   Column 271   Coefficient 48.65917969
   "001100001011000100", -- Line 1   Column 272   Coefficient 48.69140625
   "001100001011100101", -- Line 1   Column 273   Coefficient 48.72363281
   "001100001100000101", -- Line 1   Column 274   Coefficient 48.75488281
   "001100001100100110", -- Line 1   Column 275   Coefficient 48.78710938
   "001100001101000110", -- Line 1   Column 276   Coefficient 48.81835938
   "001100001101100110", -- Line 1   Column 277   Coefficient 48.84960938
   "001100001110000110", -- Line 1   Column 278   Coefficient 48.88085938
   "001100001110100110", -- Line 1   Column 279   Coefficient 48.91210938
   "001100001111000110", -- Line 1   Column 280   Coefficient 48.94335938
   "001100001111100110", -- Line 1   Column 281   Coefficient 48.97460938
   "001100010000000101", -- Line 1   Column 282   Coefficient 49.00488281
   "001100010000100101", -- Line 1   Column 283   Coefficient 49.03613281
   "001100010001000100", -- Line 1   Column 284   Coefficient 49.06640625
   "001100010001100011", -- Line 1   Column 285   Coefficient 49.09667969
   "001100010010000010", -- Line 1   Column 286   Coefficient 49.12695313
   "001100010010100001", -- Line 1   Column 287   Coefficient 49.15722656
   "001100010011000000", -- Line 1   Column 288   Coefficient 49.18750000
   "001100010011011111", -- Line 1   Column 289   Coefficient 49.21777344
   "001100010011111110", -- Line 1   Column 290   Coefficient 49.24804688
   "001100010100011101", -- Line 1   Column 291   Coefficient 49.27832031
   "001100010100111011", -- Line 1   Column 292   Coefficient 49.30761719
   "001100010101011001", -- Line 1   Column 293   Coefficient 49.33691406
   "001100010101111000", -- Line 1   Column 294   Coefficient 49.36718750
   "001100010110010110", -- Line 1   Column 295   Coefficient 49.39648438
   "001100010110110100", -- Line 1   Column 296   Coefficient 49.42578125
   "001100010111010010", -- Line 1   Column 297   Coefficient 49.45507813
   "001100010111110000", -- Line 1   Column 298   Coefficient 49.48437500
   "001100011000001110", -- Line 1   Column 299   Coefficient 49.51367188
   "001100011000101011", -- Line 1   Column 300   Coefficient 49.54199219
   "001100011001001001", -- Line 1   Column 301   Coefficient 49.57128906
   "001100011001100111", -- Line 1   Column 302   Coefficient 49.60058594
   "001100011010000100", -- Line 1   Column 303   Coefficient 49.62890625
   "001100011010100001", -- Line 1   Column 304   Coefficient 49.65722656
   "001100011010111110", -- Line 1   Column 305   Coefficient 49.68554688
   "001100011011011100", -- Line 1   Column 306   Coefficient 49.71484375
   "001100011011111001", -- Line 1   Column 307   Coefficient 49.74316406
   "001100011100010110", -- Line 1   Column 308   Coefficient 49.77148438
   "001100011100110010", -- Line 1   Column 309   Coefficient 49.79882813
   "001100011101001111", -- Line 1   Column 310   Coefficient 49.82714844
   "001100011101101100", -- Line 1   Column 311   Coefficient 49.85546875
   "001100011110001000", -- Line 1   Column 312   Coefficient 49.88281250
   "001100011110100101", -- Line 1   Column 313   Coefficient 49.91113281
   "001100011111000001", -- Line 1   Column 314   Coefficient 49.93847656
   "001100011111011101", -- Line 1   Column 315   Coefficient 49.96582031
   "001100011111111010", -- Line 1   Column 316   Coefficient 49.99414063
   "001100100000010110", -- Line 1   Column 317   Coefficient 50.02148438
   "001100100000110010", -- Line 1   Column 318   Coefficient 50.04882813
   "001100100001001110", -- Line 1   Column 319   Coefficient 50.07617188
   "001100100001101001", -- Line 1   Column 320   Coefficient 50.10253906
   "001100100010000101", -- Line 1   Column 321   Coefficient 50.12988281
   "001100100010100001", -- Line 1   Column 322   Coefficient 50.15722656
   "001100100010111100", -- Line 1   Column 323   Coefficient 50.18359375
   "001100100011011000", -- Line 1   Column 324   Coefficient 50.21093750
   "001100100011110011", -- Line 1   Column 325   Coefficient 50.23730469
   "001100100100001111", -- Line 1   Column 326   Coefficient 50.26464844
   "001100100100101010", -- Line 1   Column 327   Coefficient 50.29101563
   "001100100101000101", -- Line 1   Column 328   Coefficient 50.31738281
   "001100100101100000", -- Line 1   Column 329   Coefficient 50.34375000
   "001100100101111011", -- Line 1   Column 330   Coefficient 50.37011719
   "001100100110010110", -- Line 1   Column 331   Coefficient 50.39648438
   "001100100110110001", -- Line 1   Column 332   Coefficient 50.42285156
   "001100100111001100", -- Line 1   Column 333   Coefficient 50.44921875
   "001100100111100110", -- Line 1   Column 334   Coefficient 50.47460938
   "001100101000000001", -- Line 1   Column 335   Coefficient 50.50097656
   "001100101000011011", -- Line 1   Column 336   Coefficient 50.52636719
   "001100101000110110", -- Line 1   Column 337   Coefficient 50.55273438
   "001100101001010000", -- Line 1   Column 338   Coefficient 50.57812500
   "001100101001101010", -- Line 1   Column 339   Coefficient 50.60351563
   "001100101010000101", -- Line 1   Column 340   Coefficient 50.62988281
   "001100101010011111", -- Line 1   Column 341   Coefficient 50.65527344
   "001100101010111001", -- Line 1   Column 342   Coefficient 50.68066406
   "001100101011010011", -- Line 1   Column 343   Coefficient 50.70605469
   "001100101011101101", -- Line 1   Column 344   Coefficient 50.73144531
   "001100101100000111", -- Line 1   Column 345   Coefficient 50.75683594
   "001100101100100000", -- Line 1   Column 346   Coefficient 50.78125000
   "001100101100111010", -- Line 1   Column 347   Coefficient 50.80664063
   "001100101101010100", -- Line 1   Column 348   Coefficient 50.83203125
   "001100101101101101", -- Line 1   Column 349   Coefficient 50.85644531
   "001100101110000111", -- Line 1   Column 350   Coefficient 50.88183594
   "001100101110100000", -- Line 1   Column 351   Coefficient 50.90625000
   "001100101110111001", -- Line 1   Column 352   Coefficient 50.93066406
   "001100101111010010", -- Line 1   Column 353   Coefficient 50.95507813
   "001100101111101100", -- Line 1   Column 354   Coefficient 50.98046875
   "001100110000000101", -- Line 1   Column 355   Coefficient 51.00488281
   "001100110000011110", -- Line 1   Column 356   Coefficient 51.02929688
   "001100110000110111", -- Line 1   Column 357   Coefficient 51.05371094
   "001100110001010000", -- Line 1   Column 358   Coefficient 51.07812500
   "001100110001101000", -- Line 1   Column 359   Coefficient 51.10156250
   "001100110010000001", -- Line 1   Column 360   Coefficient 51.12597656
   "001100110010011010", -- Line 1   Column 361   Coefficient 51.15039063
   "001100110010110010", -- Line 1   Column 362   Coefficient 51.17382813
   "001100110011001011", -- Line 1   Column 363   Coefficient 51.19824219
   "001100110011100011", -- Line 1   Column 364   Coefficient 51.22167969
   "001100110011111100", -- Line 1   Column 365   Coefficient 51.24609375
   "001100110100010100", -- Line 1   Column 366   Coefficient 51.26953125
   "001100110100101100", -- Line 1   Column 367   Coefficient 51.29296875
   "001100110101000101", -- Line 1   Column 368   Coefficient 51.31738281
   "001100110101011101", -- Line 1   Column 369   Coefficient 51.34082031
   "001100110101110101", -- Line 1   Column 370   Coefficient 51.36425781
   "001100110110001101", -- Line 1   Column 371   Coefficient 51.38769531
   "001100110110100101", -- Line 1   Column 372   Coefficient 51.41113281
   "001100110110111101", -- Line 1   Column 373   Coefficient 51.43457031
   "001100110111010100", -- Line 1   Column 374   Coefficient 51.45703125
   "001100110111101100", -- Line 1   Column 375   Coefficient 51.48046875
   "001100111000000100", -- Line 1   Column 376   Coefficient 51.50390625
   "001100111000011011", -- Line 1   Column 377   Coefficient 51.52636719
   "001100111000110011", -- Line 1   Column 378   Coefficient 51.54980469
   "001100111001001011", -- Line 1   Column 379   Coefficient 51.57324219
   "001100111001100010", -- Line 1   Column 380   Coefficient 51.59570313
   "001100111001111001", -- Line 1   Column 381   Coefficient 51.61816406
   "001100111010010001", -- Line 1   Column 382   Coefficient 51.64160156
   "001100111010101000", -- Line 1   Column 383   Coefficient 51.66406250
   "001100111010111111", -- Line 1   Column 384   Coefficient 51.68652344
   "001100111011010110", -- Line 1   Column 385   Coefficient 51.70898438
   "001100111011101101", -- Line 1   Column 386   Coefficient 51.73144531
   "001100111100000100", -- Line 1   Column 387   Coefficient 51.75390625
   "001100111100011011", -- Line 1   Column 388   Coefficient 51.77636719
   "001100111100110010", -- Line 1   Column 389   Coefficient 51.79882813
   "001100111101001001", -- Line 1   Column 390   Coefficient 51.82128906
   "001100111101100000", -- Line 1   Column 391   Coefficient 51.84375000
   "001100111101110110", -- Line 1   Column 392   Coefficient 51.86523438
   "001100111110001101", -- Line 1   Column 393   Coefficient 51.88769531
   "001100111110100100", -- Line 1   Column 394   Coefficient 51.91015625
   "001100111110111010", -- Line 1   Column 395   Coefficient 51.93164063
   "001100111111010001", -- Line 1   Column 396   Coefficient 51.95410156
   "001100111111100111", -- Line 1   Column 397   Coefficient 51.97558594
   "001100111111111110", -- Line 1   Column 398   Coefficient 51.99804688
   "001101000000010100", -- Line 1   Column 399   Coefficient 52.01953125
   "001101000000101010", -- Line 1   Column 400   Coefficient 52.04101563
   "001101000001000000", -- Line 1   Column 401   Coefficient 52.06250000
   "001101000001010111", -- Line 1   Column 402   Coefficient 52.08496094
   "001101000001101101", -- Line 1   Column 403   Coefficient 52.10644531
   "001101000010000011", -- Line 1   Column 404   Coefficient 52.12792969
   "001101000010011001", -- Line 1   Column 405   Coefficient 52.14941406
   "001101000010101111", -- Line 1   Column 406   Coefficient 52.17089844
   "001101000011000100", -- Line 1   Column 407   Coefficient 52.19140625
   "001101000011011010", -- Line 1   Column 408   Coefficient 52.21289063
   "001101000011110000", -- Line 1   Column 409   Coefficient 52.23437500
   "001101000100000110", -- Line 1   Column 410   Coefficient 52.25585938
   "001101000100011011", -- Line 1   Column 411   Coefficient 52.27636719
   "001101000100110001", -- Line 1   Column 412   Coefficient 52.29785156
   "001101000101000111", -- Line 1   Column 413   Coefficient 52.31933594
   "001101000101011100", -- Line 1   Column 414   Coefficient 52.33984375
   "001101000101110010", -- Line 1   Column 415   Coefficient 52.36132813
   "001101000110000111", -- Line 1   Column 416   Coefficient 52.38183594
   "001101000110011100", -- Line 1   Column 417   Coefficient 52.40234375
   "001101000110110010", -- Line 1   Column 418   Coefficient 52.42382813
   "001101000111000111", -- Line 1   Column 419   Coefficient 52.44433594
   "001101000111011100", -- Line 1   Column 420   Coefficient 52.46484375
   "001101000111110001", -- Line 1   Column 421   Coefficient 52.48535156
   "001101001000000110", -- Line 1   Column 422   Coefficient 52.50585938
   "001101001000011011", -- Line 1   Column 423   Coefficient 52.52636719
   "001101001000110000", -- Line 1   Column 424   Coefficient 52.54687500
   "001101001001000101", -- Line 1   Column 425   Coefficient 52.56738281
   "001101001001011010", -- Line 1   Column 426   Coefficient 52.58789063
   "001101001001101111", -- Line 1   Column 427   Coefficient 52.60839844
   "001101001010000100", -- Line 1   Column 428   Coefficient 52.62890625
   "001101001010011001", -- Line 1   Column 429   Coefficient 52.64941406
   "001101001010101101", -- Line 1   Column 430   Coefficient 52.66894531
   "001101001011000010", -- Line 1   Column 431   Coefficient 52.68945313
   "001101001011010111", -- Line 1   Column 432   Coefficient 52.70996094
   "001101001011101011", -- Line 1   Column 433   Coefficient 52.72949219
   "001101001100000000", -- Line 1   Column 434   Coefficient 52.75000000
   "001101001100010100", -- Line 1   Column 435   Coefficient 52.76953125
   "001101001100101001", -- Line 1   Column 436   Coefficient 52.79003906
   "001101001100111101", -- Line 1   Column 437   Coefficient 52.80957031
   "001101001101010001", -- Line 1   Column 438   Coefficient 52.82910156
   "001101001101100110", -- Line 1   Column 439   Coefficient 52.84960938
   "001101001101111010", -- Line 1   Column 440   Coefficient 52.86914063
   "001101001110001110", -- Line 1   Column 441   Coefficient 52.88867188
   "001101001110100010", -- Line 1   Column 442   Coefficient 52.90820313
   "001101001110110110", -- Line 1   Column 443   Coefficient 52.92773438
   "001101001111001010", -- Line 1   Column 444   Coefficient 52.94726563
   "001101001111011110", -- Line 1   Column 445   Coefficient 52.96679688
   "001101001111110010", -- Line 1   Column 446   Coefficient 52.98632813
   "001101010000000110", -- Line 1   Column 447   Coefficient 53.00585938
   "001101010000011010", -- Line 1   Column 448   Coefficient 53.02539063
   "001101010000101110", -- Line 1   Column 449   Coefficient 53.04492188
   "001101010001000010", -- Line 1   Column 450   Coefficient 53.06445313
   "001101010001010110", -- Line 1   Column 451   Coefficient 53.08398438
   "001101010001101001", -- Line 1   Column 452   Coefficient 53.10253906
   "001101010001111101", -- Line 1   Column 453   Coefficient 53.12207031
   "001101010010010001", -- Line 1   Column 454   Coefficient 53.14160156
   "001101010010100100", -- Line 1   Column 455   Coefficient 53.16015625
   "001101010010111000", -- Line 1   Column 456   Coefficient 53.17968750
   "001101010011001011", -- Line 1   Column 457   Coefficient 53.19824219
   "001101010011011111", -- Line 1   Column 458   Coefficient 53.21777344
   "001101010011110010", -- Line 1   Column 459   Coefficient 53.23632813
   "001101010100000101", -- Line 1   Column 460   Coefficient 53.25488281
   "001101010100011001", -- Line 1   Column 461   Coefficient 53.27441406
   "001101010100101100", -- Line 1   Column 462   Coefficient 53.29296875
   "001101010100111111", -- Line 1   Column 463   Coefficient 53.31152344
   "001101010101010010", -- Line 1   Column 464   Coefficient 53.33007813
   "001101010101100101", -- Line 1   Column 465   Coefficient 53.34863281
   "001101010101111001", -- Line 1   Column 466   Coefficient 53.36816406
   "001101010110001100", -- Line 1   Column 467   Coefficient 53.38671875
   "001101010110011111", -- Line 1   Column 468   Coefficient 53.40527344
   "001101010110110010", -- Line 1   Column 469   Coefficient 53.42382813
   "001101010111000101", -- Line 1   Column 470   Coefficient 53.44238281
   "001101010111010111", -- Line 1   Column 471   Coefficient 53.45996094
   "001101010111101010", -- Line 1   Column 472   Coefficient 53.47851563
   "001101010111111101", -- Line 1   Column 473   Coefficient 53.49707031
   "001101011000010000", -- Line 1   Column 474   Coefficient 53.51562500
   "001101011000100011", -- Line 1   Column 475   Coefficient 53.53417969
   "001101011000110101", -- Line 1   Column 476   Coefficient 53.55175781
   "001101011001001000", -- Line 1   Column 477   Coefficient 53.57031250
   "001101011001011011", -- Line 1   Column 478   Coefficient 53.58886719
   "001101011001101101", -- Line 1   Column 479   Coefficient 53.60644531
   "001101011010000000", -- Line 1   Column 480   Coefficient 53.62500000
   "001101011010010010", -- Line 1   Column 481   Coefficient 53.64257813
   "001101011010100101", -- Line 1   Column 482   Coefficient 53.66113281
   "001101011010110111", -- Line 1   Column 483   Coefficient 53.67871094
   "001101011011001010", -- Line 1   Column 484   Coefficient 53.69726563
   "001101011011011100", -- Line 1   Column 485   Coefficient 53.71484375
   "001101011011101110", -- Line 1   Column 486   Coefficient 53.73242188
   "001101011100000001", -- Line 1   Column 487   Coefficient 53.75097656
   "001101011100010011", -- Line 1   Column 488   Coefficient 53.76855469
   "001101011100100101", -- Line 1   Column 489   Coefficient 53.78613281
   "001101011100110111", -- Line 1   Column 490   Coefficient 53.80371094
   "001101011101001001", -- Line 1   Column 491   Coefficient 53.82128906
   "001101011101011011", -- Line 1   Column 492   Coefficient 53.83886719
   "001101011101101110", -- Line 1   Column 493   Coefficient 53.85742188
   "001101011110000000", -- Line 1   Column 494   Coefficient 53.87500000
   "001101011110010010", -- Line 1   Column 495   Coefficient 53.89257813
   "001101011110100011", -- Line 1   Column 496   Coefficient 53.90917969
   "001101011110110101", -- Line 1   Column 497   Coefficient 53.92675781
   "001101011111000111", -- Line 1   Column 498   Coefficient 53.94433594
   "001101011111011001", -- Line 1   Column 499   Coefficient 53.96191406
   "001101011111101011", -- Line 1   Column 500   Coefficient 53.97949219
   "001101011111111101", -- Line 1   Column 501   Coefficient 53.99707031
   "001101100000001110", -- Line 1   Column 502   Coefficient 54.01367188
   "001101100000100000", -- Line 1   Column 503   Coefficient 54.03125000
   "001101100000110010", -- Line 1   Column 504   Coefficient 54.04882813
   "001101100001000011", -- Line 1   Column 505   Coefficient 54.06542969
   "001101100001010101", -- Line 1   Column 506   Coefficient 54.08300781
   "001101100001100111", -- Line 1   Column 507   Coefficient 54.10058594
   "001101100001111000", -- Line 1   Column 508   Coefficient 54.11718750
   "001101100010001010", -- Line 1   Column 509   Coefficient 54.13476563
   "001101100010011011", -- Line 1   Column 510   Coefficient 54.15136719
   "001101100010101100", -- Line 1   Column 511   Coefficient 54.16796875
   "001101100010111110", -- Line 1   Column 512   Coefficient 54.18554688
   "001101100011001111", -- Line 1   Column 513   Coefficient 54.20214844
   "001101100011100001", -- Line 1   Column 514   Coefficient 54.21972656
   "001101100011110010", -- Line 1   Column 515   Coefficient 54.23632813
   "001101100100000011", -- Line 1   Column 516   Coefficient 54.25292969
   "001101100100010100", -- Line 1   Column 517   Coefficient 54.26953125
   "001101100100100101", -- Line 1   Column 518   Coefficient 54.28613281
   "001101100100110111", -- Line 1   Column 519   Coefficient 54.30371094
   "001101100101001000", -- Line 1   Column 520   Coefficient 54.32031250
   "001101100101011001", -- Line 1   Column 521   Coefficient 54.33691406
   "001101100101101010", -- Line 1   Column 522   Coefficient 54.35351563
   "001101100101111011", -- Line 1   Column 523   Coefficient 54.37011719
   "001101100110001100", -- Line 1   Column 524   Coefficient 54.38671875
   "001101100110011101", -- Line 1   Column 525   Coefficient 54.40332031
   "001101100110101110", -- Line 1   Column 526   Coefficient 54.41992188
   "001101100110111111", -- Line 1   Column 527   Coefficient 54.43652344
   "001101100111010000", -- Line 1   Column 528   Coefficient 54.45312500
   "001101100111100000", -- Line 1   Column 529   Coefficient 54.46875000
   "001101100111110001", -- Line 1   Column 530   Coefficient 54.48535156
   "001101101000000010", -- Line 1   Column 531   Coefficient 54.50195313
   "001101101000010011", -- Line 1   Column 532   Coefficient 54.51855469
   "001101101000100011", -- Line 1   Column 533   Coefficient 54.53417969
   "001101101000110100", -- Line 1   Column 534   Coefficient 54.55078125
   "001101101001000101", -- Line 1   Column 535   Coefficient 54.56738281
   "001101101001010101", -- Line 1   Column 536   Coefficient 54.58300781
   "001101101001100110", -- Line 1   Column 537   Coefficient 54.59960938
   "001101101001110110", -- Line 1   Column 538   Coefficient 54.61523438
   "001101101010000111", -- Line 1   Column 539   Coefficient 54.63183594
   "001101101010010111", -- Line 1   Column 540   Coefficient 54.64746094
   "001101101010101000", -- Line 1   Column 541   Coefficient 54.66406250
   "001101101010111000", -- Line 1   Column 542   Coefficient 54.67968750
   "001101101011001001", -- Line 1   Column 543   Coefficient 54.69628906
   "001101101011011001", -- Line 1   Column 544   Coefficient 54.71191406
   "001101101011101001", -- Line 1   Column 545   Coefficient 54.72753906
   "001101101011111010", -- Line 1   Column 546   Coefficient 54.74414063
   "001101101100001010", -- Line 1   Column 547   Coefficient 54.75976563
   "001101101100011010", -- Line 1   Column 548   Coefficient 54.77539063
   "001101101100101010", -- Line 1   Column 549   Coefficient 54.79101563
   "001101101100111011", -- Line 1   Column 550   Coefficient 54.80761719
   "001101101101001011", -- Line 1   Column 551   Coefficient 54.82324219
   "001101101101011011", -- Line 1   Column 552   Coefficient 54.83886719
   "001101101101101011", -- Line 1   Column 553   Coefficient 54.85449219
   "001101101101111011", -- Line 1   Column 554   Coefficient 54.87011719
   "001101101110001011", -- Line 1   Column 555   Coefficient 54.88574219
   "001101101110011011", -- Line 1   Column 556   Coefficient 54.90136719
   "001101101110101011", -- Line 1   Column 557   Coefficient 54.91699219
   "001101101110111011", -- Line 1   Column 558   Coefficient 54.93261719
   "001101101111001011", -- Line 1   Column 559   Coefficient 54.94824219
   "001101101111011011", -- Line 1   Column 560   Coefficient 54.96386719
   "001101101111101011", -- Line 1   Column 561   Coefficient 54.97949219
   "001101101111111011", -- Line 1   Column 562   Coefficient 54.99511719
   "001101110000001010", -- Line 1   Column 563   Coefficient 55.00976563
   "001101110000011010", -- Line 1   Column 564   Coefficient 55.02539063
   "001101110000101010", -- Line 1   Column 565   Coefficient 55.04101563
   "001101110000111010", -- Line 1   Column 566   Coefficient 55.05664063
   "001101110001001001", -- Line 1   Column 567   Coefficient 55.07128906
   "001101110001011001", -- Line 1   Column 568   Coefficient 55.08691406
   "001101110001101001", -- Line 1   Column 569   Coefficient 55.10253906
   "001101110001111000", -- Line 1   Column 570   Coefficient 55.11718750
   "001101110010001000", -- Line 1   Column 571   Coefficient 55.13281250
   "001101110010010111", -- Line 1   Column 572   Coefficient 55.14746094
   "001101110010100111", -- Line 1   Column 573   Coefficient 55.16308594
   "001101110010110111", -- Line 1   Column 574   Coefficient 55.17871094
   "001101110011000110", -- Line 1   Column 575   Coefficient 55.19335938
   "001101110011010101", -- Line 1   Column 576   Coefficient 55.20800781
   "001101110011100101", -- Line 1   Column 577   Coefficient 55.22363281
   "001101110011110100", -- Line 1   Column 578   Coefficient 55.23828125
   "001101110100000100", -- Line 1   Column 579   Coefficient 55.25390625
   "001101110100010011", -- Line 1   Column 580   Coefficient 55.26855469
   "001101110100100010", -- Line 1   Column 581   Coefficient 55.28320313
   "001101110100110010", -- Line 1   Column 582   Coefficient 55.29882813
   "001101110101000001", -- Line 1   Column 583   Coefficient 55.31347656
   "001101110101010000", -- Line 1   Column 584   Coefficient 55.32812500
   "001101110101011111", -- Line 1   Column 585   Coefficient 55.34277344
   "001101110101101111", -- Line 1   Column 586   Coefficient 55.35839844
   "001101110101111110", -- Line 1   Column 587   Coefficient 55.37304688
   "001101110110001101", -- Line 1   Column 588   Coefficient 55.38769531
   "001101110110011100", -- Line 1   Column 589   Coefficient 55.40234375
   "001101110110101011", -- Line 1   Column 590   Coefficient 55.41699219
   "001101110110111010", -- Line 1   Column 591   Coefficient 55.43164063
   "001101110111001001", -- Line 1   Column 592   Coefficient 55.44628906
   "001101110111011000", -- Line 1   Column 593   Coefficient 55.46093750
   "001101110111100111", -- Line 1   Column 594   Coefficient 55.47558594
   "001101110111110110", -- Line 1   Column 595   Coefficient 55.49023438
   "001101111000000101", -- Line 1   Column 596   Coefficient 55.50488281
   "001101111000010100", -- Line 1   Column 597   Coefficient 55.51953125
   "001101111000100011", -- Line 1   Column 598   Coefficient 55.53417969
   "001101111000110010", -- Line 1   Column 599   Coefficient 55.54882813
   "001101111001000001", -- Line 1   Column 600   Coefficient 55.56347656
   "001101111001001111", -- Line 1   Column 601   Coefficient 55.57714844
   "001101111001011110", -- Line 1   Column 602   Coefficient 55.59179688
   "001101111001101101", -- Line 1   Column 603   Coefficient 55.60644531
   "001101111001111100", -- Line 1   Column 604   Coefficient 55.62109375
   "001101111010001010", -- Line 1   Column 605   Coefficient 55.63476563
   "001101111010011001", -- Line 1   Column 606   Coefficient 55.64941406
   "001101111010101000", -- Line 1   Column 607   Coefficient 55.66406250
   "001101111010110110", -- Line 1   Column 608   Coefficient 55.67773438
   "001101111011000101", -- Line 1   Column 609   Coefficient 55.69238281
   "001101111011010100", -- Line 1   Column 610   Coefficient 55.70703125
   "001101111011100010", -- Line 1   Column 611   Coefficient 55.72070313
   "001101111011110001", -- Line 1   Column 612   Coefficient 55.73535156
   "001101111011111111", -- Line 1   Column 613   Coefficient 55.74902344
   "001101111100001110", -- Line 1   Column 614   Coefficient 55.76367188
   "001101111100011100", -- Line 1   Column 615   Coefficient 55.77734375
   "001101111100101011", -- Line 1   Column 616   Coefficient 55.79199219
   "001101111100111001", -- Line 1   Column 617   Coefficient 55.80566406
   "001101111101000111", -- Line 1   Column 618   Coefficient 55.81933594
   "001101111101010110", -- Line 1   Column 619   Coefficient 55.83398438
   "001101111101100100", -- Line 1   Column 620   Coefficient 55.84765625
   "001101111101110011", -- Line 1   Column 621   Coefficient 55.86230469
   "001101111110000001", -- Line 1   Column 622   Coefficient 55.87597656
   "001101111110001111", -- Line 1   Column 623   Coefficient 55.88964844
   "001101111110011101", -- Line 1   Column 624   Coefficient 55.90332031
   "001101111110101100", -- Line 1   Column 625   Coefficient 55.91796875
   "001101111110111010", -- Line 1   Column 626   Coefficient 55.93164063
   "001101111111001000", -- Line 1   Column 627   Coefficient 55.94531250
   "001101111111010110", -- Line 1   Column 628   Coefficient 55.95898438
   "001101111111100100", -- Line 1   Column 629   Coefficient 55.97265625
   "001101111111110010", -- Line 1   Column 630   Coefficient 55.98632813
   "001110000000000001", -- Line 1   Column 631   Coefficient 56.00097656
   "001110000000001111", -- Line 1   Column 632   Coefficient 56.01464844
   "001110000000011101", -- Line 1   Column 633   Coefficient 56.02832031
   "001110000000101011", -- Line 1   Column 634   Coefficient 56.04199219
   "001110000000111001", -- Line 1   Column 635   Coefficient 56.05566406
   "001110000001000111", -- Line 1   Column 636   Coefficient 56.06933594
   "001110000001010101", -- Line 1   Column 637   Coefficient 56.08300781
   "001110000001100011", -- Line 1   Column 638   Coefficient 56.09667969
   "001110000001110001", -- Line 1   Column 639   Coefficient 56.11035156
   "001110000001111111", -- Line 1   Column 640   Coefficient 56.12402344
   "001110000010001100", -- Line 1   Column 641   Coefficient 56.13671875
   "001110000010011010", -- Line 1   Column 642   Coefficient 56.15039063
   "001110000010101000", -- Line 1   Column 643   Coefficient 56.16406250
   "001110000010110110", -- Line 1   Column 644   Coefficient 56.17773438
   "001110000011000100", -- Line 1   Column 645   Coefficient 56.19140625
   "001110000011010010", -- Line 1   Column 646   Coefficient 56.20507813
   "001110000011011111", -- Line 1   Column 647   Coefficient 56.21777344
   "001110000011101101", -- Line 1   Column 648   Coefficient 56.23144531
   "001110000011111011", -- Line 1   Column 649   Coefficient 56.24511719
   "001110000100001000", -- Line 1   Column 650   Coefficient 56.25781250
   "001110000100010110", -- Line 1   Column 651   Coefficient 56.27148438
   "001110000100100100", -- Line 1   Column 652   Coefficient 56.28515625
   "001110000100110001", -- Line 1   Column 653   Coefficient 56.29785156
   "001110000100111111", -- Line 1   Column 654   Coefficient 56.31152344
   "001110000101001101", -- Line 1   Column 655   Coefficient 56.32519531
   "001110000101011010", -- Line 1   Column 656   Coefficient 56.33789063
   "001110000101101000", -- Line 1   Column 657   Coefficient 56.35156250
   "001110000101110101", -- Line 1   Column 658   Coefficient 56.36425781
   "001110000110000011", -- Line 1   Column 659   Coefficient 56.37792969
   "001110000110010000", -- Line 1   Column 660   Coefficient 56.39062500
   "001110000110011110", -- Line 1   Column 661   Coefficient 56.40429688
   "001110000110101011", -- Line 1   Column 662   Coefficient 56.41699219
   "001110000110111001", -- Line 1   Column 663   Coefficient 56.43066406
   "001110000111000110", -- Line 1   Column 664   Coefficient 56.44335938
   "001110000111010011", -- Line 1   Column 665   Coefficient 56.45605469
   "001110000111100001", -- Line 1   Column 666   Coefficient 56.46972656
   "001110000111101110", -- Line 1   Column 667   Coefficient 56.48242188
   "001110000111111011", -- Line 1   Column 668   Coefficient 56.49511719
   "001110001000001001", -- Line 1   Column 669   Coefficient 56.50878906
   "001110001000010110", -- Line 1   Column 670   Coefficient 56.52148438
   "001110001000100011", -- Line 1   Column 671   Coefficient 56.53417969
   "001110001000110001", -- Line 1   Column 672   Coefficient 56.54785156
   "001110001000111110", -- Line 1   Column 673   Coefficient 56.56054688
   "001110001001001011", -- Line 1   Column 674   Coefficient 56.57324219
   "001110001001011000", -- Line 1   Column 675   Coefficient 56.58593750
   "001110001001100101", -- Line 1   Column 676   Coefficient 56.59863281
   "001110001001110010", -- Line 1   Column 677   Coefficient 56.61132813
   "001110001010000000", -- Line 1   Column 678   Coefficient 56.62500000
   "001110001010001101", -- Line 1   Column 679   Coefficient 56.63769531
   "001110001010011010", -- Line 1   Column 680   Coefficient 56.65039063
   "001110001010100111", -- Line 1   Column 681   Coefficient 56.66308594
   "001110001010110100", -- Line 1   Column 682   Coefficient 56.67578125
   "001110001011000001", -- Line 1   Column 683   Coefficient 56.68847656
   "001110001011001110", -- Line 1   Column 684   Coefficient 56.70117188
   "001110001011011011", -- Line 1   Column 685   Coefficient 56.71386719
   "001110001011101000", -- Line 1   Column 686   Coefficient 56.72656250
   "001110001011110101", -- Line 1   Column 687   Coefficient 56.73925781
   "001110001100000010", -- Line 1   Column 688   Coefficient 56.75195313
   "001110001100001111", -- Line 1   Column 689   Coefficient 56.76464844
   "001110001100011100", -- Line 1   Column 690   Coefficient 56.77734375
   "001110001100101001", -- Line 1   Column 691   Coefficient 56.79003906
   "001110001100110101", -- Line 1   Column 692   Coefficient 56.80175781
   "001110001101000010", -- Line 1   Column 693   Coefficient 56.81445313
   "001110001101001111", -- Line 1   Column 694   Coefficient 56.82714844
   "001110001101011100", -- Line 1   Column 695   Coefficient 56.83984375
   "001110001101101001", -- Line 1   Column 696   Coefficient 56.85253906
   "001110001101110101", -- Line 1   Column 697   Coefficient 56.86425781
   "001110001110000010", -- Line 1   Column 698   Coefficient 56.87695313
   "001110001110001111", -- Line 1   Column 699   Coefficient 56.88964844
   "001110001110011100", -- Line 1   Column 700   Coefficient 56.90234375
   "001110001110101000", -- Line 1   Column 701   Coefficient 56.91406250
   "001110001110110101", -- Line 1   Column 702   Coefficient 56.92675781
   "001110001111000010", -- Line 1   Column 703   Coefficient 56.93945313
   "001110001111001110", -- Line 1   Column 704   Coefficient 56.95117188
   "001110001111011011", -- Line 1   Column 705   Coefficient 56.96386719
   "001110001111101000", -- Line 1   Column 706   Coefficient 56.97656250
   "001110001111110100", -- Line 1   Column 707   Coefficient 56.98828125
   "001110010000000001", -- Line 1   Column 708   Coefficient 57.00097656
   "001110010000001101", -- Line 1   Column 709   Coefficient 57.01269531
   "001110010000011010", -- Line 1   Column 710   Coefficient 57.02539063
   "001110010000100110", -- Line 1   Column 711   Coefficient 57.03710938
   "001110010000110011", -- Line 1   Column 712   Coefficient 57.04980469
   "001110010000111111", -- Line 1   Column 713   Coefficient 57.06152344
   "001110010001001100", -- Line 1   Column 714   Coefficient 57.07421875
   "001110010001011000", -- Line 1   Column 715   Coefficient 57.08593750
   "001110010001100101", -- Line 1   Column 716   Coefficient 57.09863281
   "001110010001110001", -- Line 1   Column 717   Coefficient 57.11035156
   "001110010001111101", -- Line 1   Column 718   Coefficient 57.12207031
   "001110010010001010", -- Line 1   Column 719   Coefficient 57.13476563
   "001110010010010110", -- Line 1   Column 720   Coefficient 57.14648438
   "001110010010100011", -- Line 1   Column 721   Coefficient 57.15917969
   "001110010010101111", -- Line 1   Column 722   Coefficient 57.17089844
   "001110010010111011", -- Line 1   Column 723   Coefficient 57.18261719
   "001110010011000111", -- Line 1   Column 724   Coefficient 57.19433594
   "001110010011010100", -- Line 1   Column 725   Coefficient 57.20703125
   "001110010011100000", -- Line 1   Column 726   Coefficient 57.21875000
   "001110010011101100", -- Line 1   Column 727   Coefficient 57.23046875
   "001110010011111000", -- Line 1   Column 728   Coefficient 57.24218750
   "001110010100000101", -- Line 1   Column 729   Coefficient 57.25488281
   "001110010100010001", -- Line 1   Column 730   Coefficient 57.26660156
   "001110010100011101", -- Line 1   Column 731   Coefficient 57.27832031
   "001110010100101001", -- Line 1   Column 732   Coefficient 57.29003906
   "001110010100110101", -- Line 1   Column 733   Coefficient 57.30175781
   "001110010101000001", -- Line 1   Column 734   Coefficient 57.31347656
   "001110010101001110", -- Line 1   Column 735   Coefficient 57.32617188
   "001110010101011010", -- Line 1   Column 736   Coefficient 57.33789063
   "001110010101100110", -- Line 1   Column 737   Coefficient 57.34960938
   "001110010101110010", -- Line 1   Column 738   Coefficient 57.36132813
   "001110010101111110", -- Line 1   Column 739   Coefficient 57.37304688
   "001110010110001010", -- Line 1   Column 740   Coefficient 57.38476563
   "001110010110010110", -- Line 1   Column 741   Coefficient 57.39648438
   "001110010110100010", -- Line 1   Column 742   Coefficient 57.40820313
   "001110010110101110", -- Line 1   Column 743   Coefficient 57.41992188
   "001110010110111010", -- Line 1   Column 744   Coefficient 57.43164063
   "001110010111000110", -- Line 1   Column 745   Coefficient 57.44335938
   "001110010111010010", -- Line 1   Column 746   Coefficient 57.45507813
   "001110010111011110", -- Line 1   Column 747   Coefficient 57.46679688
   "001110010111101010", -- Line 1   Column 748   Coefficient 57.47851563
   "001110010111110101", -- Line 1   Column 749   Coefficient 57.48925781
   "001110011000000001", -- Line 1   Column 750   Coefficient 57.50097656
   "001110011000001101", -- Line 1   Column 751   Coefficient 57.51269531
   "001110011000011001", -- Line 1   Column 752   Coefficient 57.52441406
   "001110011000100101", -- Line 1   Column 753   Coefficient 57.53613281
   "001110011000110001", -- Line 1   Column 754   Coefficient 57.54785156
   "001110011000111100", -- Line 1   Column 755   Coefficient 57.55859375
   "001110011001001000", -- Line 1   Column 756   Coefficient 57.57031250
   "001110011001010100", -- Line 1   Column 757   Coefficient 57.58203125
   "001110011001100000", -- Line 1   Column 758   Coefficient 57.59375000
   "001110011001101011", -- Line 1   Column 759   Coefficient 57.60449219
   "001110011001110111", -- Line 1   Column 760   Coefficient 57.61621094
   "001110011010000011", -- Line 1   Column 761   Coefficient 57.62792969
   "001110011010001110", -- Line 1   Column 762   Coefficient 57.63867188
   "001110011010011010", -- Line 1   Column 763   Coefficient 57.65039063
   "001110011010100110", -- Line 1   Column 764   Coefficient 57.66210938
   "001110011010110001", -- Line 1   Column 765   Coefficient 57.67285156
   "001110011010111101", -- Line 1   Column 766   Coefficient 57.68457031
   "001110011011001001", -- Line 1   Column 767   Coefficient 57.69628906
   "001110011011010100", -- Line 1   Column 768   Coefficient 57.70703125
   "001110011011100000", -- Line 1   Column 769   Coefficient 57.71875000
   "001110011011101011", -- Line 1   Column 770   Coefficient 57.72949219
   "001110011011110111", -- Line 1   Column 771   Coefficient 57.74121094
   "001110011100000010", -- Line 1   Column 772   Coefficient 57.75195313
   "001110011100001110", -- Line 1   Column 773   Coefficient 57.76367188
   "001110011100011001", -- Line 1   Column 774   Coefficient 57.77441406
   "001110011100100101", -- Line 1   Column 775   Coefficient 57.78613281
   "001110011100110000", -- Line 1   Column 776   Coefficient 57.79687500
   "001110011100111100", -- Line 1   Column 777   Coefficient 57.80859375
   "001110011101000111", -- Line 1   Column 778   Coefficient 57.81933594
   "001110011101010011", -- Line 1   Column 779   Coefficient 57.83105469
   "001110011101011110", -- Line 1   Column 780   Coefficient 57.84179688
   "001110011101101001", -- Line 1   Column 781   Coefficient 57.85253906
   "001110011101110101", -- Line 1   Column 782   Coefficient 57.86425781
   "001110011110000000", -- Line 1   Column 783   Coefficient 57.87500000
   "001110011110001100", -- Line 1   Column 784   Coefficient 57.88671875
   "001110011110010111", -- Line 1   Column 785   Coefficient 57.89746094
   "001110011110100010", -- Line 1   Column 786   Coefficient 57.90820313
   "001110011110101110", -- Line 1   Column 787   Coefficient 57.91992188
   "001110011110111001", -- Line 1   Column 788   Coefficient 57.93066406
   "001110011111000100", -- Line 1   Column 789   Coefficient 57.94140625
   "001110011111001111", -- Line 1   Column 790   Coefficient 57.95214844
   "001110011111011011", -- Line 1   Column 791   Coefficient 57.96386719
   "001110011111100110", -- Line 1   Column 792   Coefficient 57.97460938
   "001110011111110001", -- Line 1   Column 793   Coefficient 57.98535156
   "001110011111111100", -- Line 1   Column 794   Coefficient 57.99609375
   "001110100000001000", -- Line 1   Column 795   Coefficient 58.00781250
   "001110100000010011", -- Line 1   Column 796   Coefficient 58.01855469
   "001110100000011110", -- Line 1   Column 797   Coefficient 58.02929688
   "001110100000101001", -- Line 1   Column 798   Coefficient 58.04003906
   "001110100000110100", -- Line 1   Column 799   Coefficient 58.05078125
   "001110100000111111", -- Line 1   Column 800   Coefficient 58.06152344
   "001110100001001010", -- Line 1   Column 801   Coefficient 58.07226563
   "001110100001010101", -- Line 1   Column 802   Coefficient 58.08300781
   "001110100001100001", -- Line 1   Column 803   Coefficient 58.09472656
   "001110100001101100", -- Line 1   Column 804   Coefficient 58.10546875
   "001110100001110111", -- Line 1   Column 805   Coefficient 58.11621094
   "001110100010000010", -- Line 1   Column 806   Coefficient 58.12695313
   "001110100010001101", -- Line 1   Column 807   Coefficient 58.13769531
   "001110100010011000", -- Line 1   Column 808   Coefficient 58.14843750
   "001110100010100011", -- Line 1   Column 809   Coefficient 58.15917969
   "001110100010101110", -- Line 1   Column 810   Coefficient 58.16992188
   "001110100010111001", -- Line 1   Column 811   Coefficient 58.18066406
   "001110100011000100", -- Line 1   Column 812   Coefficient 58.19140625
   "001110100011001111", -- Line 1   Column 813   Coefficient 58.20214844
   "001110100011011010", -- Line 1   Column 814   Coefficient 58.21289063
   "001110100011100101", -- Line 1   Column 815   Coefficient 58.22363281
   "001110100011101111", -- Line 1   Column 816   Coefficient 58.23339844
   "001110100011111010", -- Line 1   Column 817   Coefficient 58.24414063
   "001110100100000101", -- Line 1   Column 818   Coefficient 58.25488281
   "001110100100010000", -- Line 1   Column 819   Coefficient 58.26562500
   "001110100100011011", -- Line 1   Column 820   Coefficient 58.27636719
   "001110100100100110", -- Line 1   Column 821   Coefficient 58.28710938
   "001110100100110001", -- Line 1   Column 822   Coefficient 58.29785156
   "001110100100111011", -- Line 1   Column 823   Coefficient 58.30761719
   "001110100101000110", -- Line 1   Column 824   Coefficient 58.31835938
   "001110100101010001", -- Line 1   Column 825   Coefficient 58.32910156
   "001110100101011100", -- Line 1   Column 826   Coefficient 58.33984375
   "001110100101100111", -- Line 1   Column 827   Coefficient 58.35058594
   "001110100101110001", -- Line 1   Column 828   Coefficient 58.36035156
   "001110100101111100", -- Line 1   Column 829   Coefficient 58.37109375
   "001110100110000111", -- Line 1   Column 830   Coefficient 58.38183594
   "001110100110010001", -- Line 1   Column 831   Coefficient 58.39160156
   "001110100110011100", -- Line 1   Column 832   Coefficient 58.40234375
   "001110100110100111", -- Line 1   Column 833   Coefficient 58.41308594
   "001110100110110001", -- Line 1   Column 834   Coefficient 58.42285156
   "001110100110111100", -- Line 1   Column 835   Coefficient 58.43359375
   "001110100111000111", -- Line 1   Column 836   Coefficient 58.44433594
   "001110100111010001", -- Line 1   Column 837   Coefficient 58.45410156
   "001110100111011100", -- Line 1   Column 838   Coefficient 58.46484375
   "001110100111100111", -- Line 1   Column 839   Coefficient 58.47558594
   "001110100111110001", -- Line 1   Column 840   Coefficient 58.48535156
   "001110100111111100", -- Line 1   Column 841   Coefficient 58.49609375
   "001110101000000110", -- Line 1   Column 842   Coefficient 58.50585938
   "001110101000010001", -- Line 1   Column 843   Coefficient 58.51660156
   "001110101000011011", -- Line 1   Column 844   Coefficient 58.52636719
   "001110101000100110", -- Line 1   Column 845   Coefficient 58.53710938
   "001110101000110001", -- Line 1   Column 846   Coefficient 58.54785156
   "001110101000111011", -- Line 1   Column 847   Coefficient 58.55761719
   "001110101001000110", -- Line 1   Column 848   Coefficient 58.56835938
   "001110101001010000", -- Line 1   Column 849   Coefficient 58.57812500
   "001110101001011010", -- Line 1   Column 850   Coefficient 58.58789063
   "001110101001100101", -- Line 1   Column 851   Coefficient 58.59863281
   "001110101001101111", -- Line 1   Column 852   Coefficient 58.60839844
   "001110101001111010", -- Line 1   Column 853   Coefficient 58.61914063
   "001110101010000100", -- Line 1   Column 854   Coefficient 58.62890625
   "001110101010001111", -- Line 1   Column 855   Coefficient 58.63964844
   "001110101010011001", -- Line 1   Column 856   Coefficient 58.64941406
   "001110101010100011", -- Line 1   Column 857   Coefficient 58.65917969
   "001110101010101110", -- Line 1   Column 858   Coefficient 58.66992188
   "001110101010111000", -- Line 1   Column 859   Coefficient 58.67968750
   "001110101011000011", -- Line 1   Column 860   Coefficient 58.69042969
   "001110101011001101", -- Line 1   Column 861   Coefficient 58.70019531
   "001110101011010111", -- Line 1   Column 862   Coefficient 58.70996094
   "001110101011100010", -- Line 1   Column 863   Coefficient 58.72070313
   "001110101011101100", -- Line 1   Column 864   Coefficient 58.73046875
   "001110101011110110", -- Line 1   Column 865   Coefficient 58.74023438
   "001110101100000000", -- Line 1   Column 866   Coefficient 58.75000000
   "001110101100001011", -- Line 1   Column 867   Coefficient 58.76074219
   "001110101100010101", -- Line 1   Column 868   Coefficient 58.77050781
   "001110101100011111", -- Line 1   Column 869   Coefficient 58.78027344
   "001110101100101001", -- Line 1   Column 870   Coefficient 58.79003906
   "001110101100110100", -- Line 1   Column 871   Coefficient 58.80078125
   "001110101100111110", -- Line 1   Column 872   Coefficient 58.81054688
   "001110101101001000", -- Line 1   Column 873   Coefficient 58.82031250
   "001110101101010010", -- Line 1   Column 874   Coefficient 58.83007813
   "001110101101011100", -- Line 1   Column 875   Coefficient 58.83984375
   "001110101101100110", -- Line 1   Column 876   Coefficient 58.84960938
   "001110101101110001", -- Line 1   Column 877   Coefficient 58.86035156
   "001110101101111011", -- Line 1   Column 878   Coefficient 58.87011719
   "001110101110000101", -- Line 1   Column 879   Coefficient 58.87988281
   "001110101110001111", -- Line 1   Column 880   Coefficient 58.88964844
   "001110101110011001", -- Line 1   Column 881   Coefficient 58.89941406
   "001110101110100011", -- Line 1   Column 882   Coefficient 58.90917969
   "001110101110101101", -- Line 1   Column 883   Coefficient 58.91894531
   "001110101110110111", -- Line 1   Column 884   Coefficient 58.92871094
   "001110101111000001", -- Line 1   Column 885   Coefficient 58.93847656
   "001110101111001011", -- Line 1   Column 886   Coefficient 58.94824219
   "001110101111010101", -- Line 1   Column 887   Coefficient 58.95800781
   "001110101111011111", -- Line 1   Column 888   Coefficient 58.96777344
   "001110101111101010", -- Line 1   Column 889   Coefficient 58.97851563
   "001110101111110100", -- Line 1   Column 890   Coefficient 58.98828125
   "001110101111111101", -- Line 1   Column 891   Coefficient 58.99707031
   "001110110000000111", -- Line 1   Column 892   Coefficient 59.00683594
   "001110110000010001", -- Line 1   Column 893   Coefficient 59.01660156
   "001110110000011011", -- Line 1   Column 894   Coefficient 59.02636719
   "001110110000100101", -- Line 1   Column 895   Coefficient 59.03613281
   "001110110000101111", -- Line 1   Column 896   Coefficient 59.04589844
   "001110110000111001", -- Line 1   Column 897   Coefficient 59.05566406
   "001110110001000011", -- Line 1   Column 898   Coefficient 59.06542969
   "001110110001001101", -- Line 1   Column 899   Coefficient 59.07519531
   "001110110001010111", -- Line 1   Column 900   Coefficient 59.08496094
   "001110110001100001", -- Line 1   Column 901   Coefficient 59.09472656
   "001110110001101011", -- Line 1   Column 902   Coefficient 59.10449219
   "001110110001110100", -- Line 1   Column 903   Coefficient 59.11328125
   "001110110001111110", -- Line 1   Column 904   Coefficient 59.12304688
   "001110110010001000", -- Line 1   Column 905   Coefficient 59.13281250
   "001110110010010010", -- Line 1   Column 906   Coefficient 59.14257813
   "001110110010011100", -- Line 1   Column 907   Coefficient 59.15234375
   "001110110010100110", -- Line 1   Column 908   Coefficient 59.16210938
   "001110110010101111", -- Line 1   Column 909   Coefficient 59.17089844
   "001110110010111001", -- Line 1   Column 910   Coefficient 59.18066406
   "001110110011000011", -- Line 1   Column 911   Coefficient 59.19042969
   "001110110011001101", -- Line 1   Column 912   Coefficient 59.20019531
   "001110110011010110", -- Line 1   Column 913   Coefficient 59.20898438
   "001110110011100000", -- Line 1   Column 914   Coefficient 59.21875000
   "001110110011101010", -- Line 1   Column 915   Coefficient 59.22851563
   "001110110011110100", -- Line 1   Column 916   Coefficient 59.23828125
   "001110110011111101", -- Line 1   Column 917   Coefficient 59.24707031
   "001110110100000111", -- Line 1   Column 918   Coefficient 59.25683594
   "001110110100010001", -- Line 1   Column 919   Coefficient 59.26660156
   "001110110100011010", -- Line 1   Column 920   Coefficient 59.27539063
   "001110110100100100", -- Line 1   Column 921   Coefficient 59.28515625
   "001110110100101110", -- Line 1   Column 922   Coefficient 59.29492188
   "001110110100110111", -- Line 1   Column 923   Coefficient 59.30371094
   "001110110101000001", -- Line 1   Column 924   Coefficient 59.31347656
   "001110110101001011", -- Line 1   Column 925   Coefficient 59.32324219
   "001110110101010100", -- Line 1   Column 926   Coefficient 59.33203125
   "001110110101011110", -- Line 1   Column 927   Coefficient 59.34179688
   "001110110101100111", -- Line 1   Column 928   Coefficient 59.35058594
   "001110110101110001", -- Line 1   Column 929   Coefficient 59.36035156
   "001110110101111011", -- Line 1   Column 930   Coefficient 59.37011719
   "001110110110000100", -- Line 1   Column 931   Coefficient 59.37890625
   "001110110110001110", -- Line 1   Column 932   Coefficient 59.38867188
   "001110110110010111", -- Line 1   Column 933   Coefficient 59.39746094
   "001110110110100001", -- Line 1   Column 934   Coefficient 59.40722656
   "001110110110101010", -- Line 1   Column 935   Coefficient 59.41601563
   "001110110110110100", -- Line 1   Column 936   Coefficient 59.42578125
   "001110110110111101", -- Line 1   Column 937   Coefficient 59.43457031
   "001110110111000111", -- Line 1   Column 938   Coefficient 59.44433594
   "001110110111010000", -- Line 1   Column 939   Coefficient 59.45312500
   "001110110111011010", -- Line 1   Column 940   Coefficient 59.46289063
   "001110110111100011", -- Line 1   Column 941   Coefficient 59.47167969
   "001110110111101101", -- Line 1   Column 942   Coefficient 59.48144531
   "001110110111110110", -- Line 1   Column 943   Coefficient 59.49023438
   "001110110111111111", -- Line 1   Column 944   Coefficient 59.49902344
   "001110111000001001", -- Line 1   Column 945   Coefficient 59.50878906
   "001110111000010010", -- Line 1   Column 946   Coefficient 59.51757813
   "001110111000011100", -- Line 1   Column 947   Coefficient 59.52734375
   "001110111000100101", -- Line 1   Column 948   Coefficient 59.53613281
   "001110111000101110", -- Line 1   Column 949   Coefficient 59.54492188
   "001110111000111000", -- Line 1   Column 950   Coefficient 59.55468750
   "001110111001000001", -- Line 1   Column 951   Coefficient 59.56347656
   "001110111001001010", -- Line 1   Column 952   Coefficient 59.57226563
   "001110111001010100", -- Line 1   Column 953   Coefficient 59.58203125
   "001110111001011101", -- Line 1   Column 954   Coefficient 59.59082031
   "001110111001100110", -- Line 1   Column 955   Coefficient 59.59960938
   "001110111001110000", -- Line 1   Column 956   Coefficient 59.60937500
   "001110111001111001", -- Line 1   Column 957   Coefficient 59.61816406
   "001110111010000010", -- Line 1   Column 958   Coefficient 59.62695313
   "001110111010001100", -- Line 1   Column 959   Coefficient 59.63671875
   "001110111010010101", -- Line 1   Column 960   Coefficient 59.64550781
   "001110111010011110", -- Line 1   Column 961   Coefficient 59.65429688
   "001110111010100111", -- Line 1   Column 962   Coefficient 59.66308594
   "001110111010110001", -- Line 1   Column 963   Coefficient 59.67285156
   "001110111010111010", -- Line 1   Column 964   Coefficient 59.68164063
   "001110111011000011", -- Line 1   Column 965   Coefficient 59.69042969
   "001110111011001100", -- Line 1   Column 966   Coefficient 59.69921875
   "001110111011010110", -- Line 1   Column 967   Coefficient 59.70898438
   "001110111011011111", -- Line 1   Column 968   Coefficient 59.71777344
   "001110111011101000", -- Line 1   Column 969   Coefficient 59.72656250
   "001110111011110001", -- Line 1   Column 970   Coefficient 59.73535156
   "001110111011111010", -- Line 1   Column 971   Coefficient 59.74414063
   "001110111100000011", -- Line 1   Column 972   Coefficient 59.75292969
   "001110111100001101", -- Line 1   Column 973   Coefficient 59.76269531
   "001110111100010110", -- Line 1   Column 974   Coefficient 59.77148438
   "001110111100011111", -- Line 1   Column 975   Coefficient 59.78027344
   "001110111100101000", -- Line 1   Column 976   Coefficient 59.78906250
   "001110111100110001", -- Line 1   Column 977   Coefficient 59.79785156
   "001110111100111010", -- Line 1   Column 978   Coefficient 59.80664063
   "001110111101000011", -- Line 1   Column 979   Coefficient 59.81542969
   "001110111101001100", -- Line 1   Column 980   Coefficient 59.82421875
   "001110111101010101", -- Line 1   Column 981   Coefficient 59.83300781
   "001110111101011110", -- Line 1   Column 982   Coefficient 59.84179688
   "001110111101100111", -- Line 1   Column 983   Coefficient 59.85058594
   "001110111101110001", -- Line 1   Column 984   Coefficient 59.86035156
   "001110111101111010", -- Line 1   Column 985   Coefficient 59.86914063
   "001110111110000011", -- Line 1   Column 986   Coefficient 59.87792969
   "001110111110001100", -- Line 1   Column 987   Coefficient 59.88671875
   "001110111110010101", -- Line 1   Column 988   Coefficient 59.89550781
   "001110111110011110", -- Line 1   Column 989   Coefficient 59.90429688
   "001110111110100111", -- Line 1   Column 990   Coefficient 59.91308594
   "001110111110110000", -- Line 1   Column 991   Coefficient 59.92187500
   "001110111110111001", -- Line 1   Column 992   Coefficient 59.93066406
   "001110111111000010", -- Line 1   Column 993   Coefficient 59.93945313
   "001110111111001010", -- Line 1   Column 994   Coefficient 59.94726563
   "001110111111010011", -- Line 1   Column 995   Coefficient 59.95605469
   "001110111111011100", -- Line 1   Column 996   Coefficient 59.96484375
   "001110111111100101", -- Line 1   Column 997   Coefficient 59.97363281
   "001110111111101110", -- Line 1   Column 998   Coefficient 59.98242188
   "001110111111110111", -- Line 1   Column 999   Coefficient 59.99121094
   "001111000000000000", -- Line 1   Column 1000   Coefficient 60.00000000
   "001111000000001001", -- Line 1   Column 1001   Coefficient 60.00878906
   "001111000000010010", -- Line 1   Column 1002   Coefficient 60.01757813
   "001111000000011011", -- Line 1   Column 1003   Coefficient 60.02636719
   "001111000000100100", -- Line 1   Column 1004   Coefficient 60.03515625
   "001111000000101100", -- Line 1   Column 1005   Coefficient 60.04296875
   "001111000000110101", -- Line 1   Column 1006   Coefficient 60.05175781
   "001111000000111110", -- Line 1   Column 1007   Coefficient 60.06054688
   "001111000001000111", -- Line 1   Column 1008   Coefficient 60.06933594
   "001111000001010000", -- Line 1   Column 1009   Coefficient 60.07812500
   "001111000001011001", -- Line 1   Column 1010   Coefficient 60.08691406
   "001111000001100001", -- Line 1   Column 1011   Coefficient 60.09472656
   "001111000001101010", -- Line 1   Column 1012   Coefficient 60.10351563
   "001111000001110011", -- Line 1   Column 1013   Coefficient 60.11230469
   "001111000001111100", -- Line 1   Column 1014   Coefficient 60.12109375
   "001111000010000100", -- Line 1   Column 1015   Coefficient 60.12890625
   "001111000010001101", -- Line 1   Column 1016   Coefficient 60.13769531
   "001111000010010110", -- Line 1   Column 1017   Coefficient 60.14648438
   "001111000010011111", -- Line 1   Column 1018   Coefficient 60.15527344
   "001111000010100111", -- Line 1   Column 1019   Coefficient 60.16308594
   "001111000010110000", -- Line 1   Column 1020   Coefficient 60.17187500
   "001111000010111001", -- Line 1   Column 1021   Coefficient 60.18066406
   "001111000011000010", -- Line 1   Column 1022   Coefficient 60.18945313
   "001111000011001010", -- Line 1   Column 1023   Coefficient 60.19726563
   "001111000011010011", -- Line 1   Column 1024   Coefficient 60.20605469
   "001111000011011100", -- Line 1   Column 1025   Coefficient 60.21484375
   "001111000011100100", -- Line 1   Column 1026   Coefficient 60.22265625
   "001111000011101101", -- Line 1   Column 1027   Coefficient 60.23144531
   "001111000011110110", -- Line 1   Column 1028   Coefficient 60.24023438
   "001111000011111110", -- Line 1   Column 1029   Coefficient 60.24804688
   "001111000100000111", -- Line 1   Column 1030   Coefficient 60.25683594
   "001111000100010000", -- Line 1   Column 1031   Coefficient 60.26562500
   "001111000100011000", -- Line 1   Column 1032   Coefficient 60.27343750
   "001111000100100001", -- Line 1   Column 1033   Coefficient 60.28222656
   "001111000100101001", -- Line 1   Column 1034   Coefficient 60.29003906
   "001111000100110010", -- Line 1   Column 1035   Coefficient 60.29882813
   "001111000100111011", -- Line 1   Column 1036   Coefficient 60.30761719
   "001111000101000011", -- Line 1   Column 1037   Coefficient 60.31542969
   "001111000101001100", -- Line 1   Column 1038   Coefficient 60.32421875
   "001111000101010100", -- Line 1   Column 1039   Coefficient 60.33203125
   "001111000101011101", -- Line 1   Column 1040   Coefficient 60.34082031
   "001111000101100101", -- Line 1   Column 1041   Coefficient 60.34863281
   "001111000101101110", -- Line 1   Column 1042   Coefficient 60.35742188
   "001111000101110110", -- Line 1   Column 1043   Coefficient 60.36523438
   "001111000101111111", -- Line 1   Column 1044   Coefficient 60.37402344
   "001111000110001000", -- Line 1   Column 1045   Coefficient 60.38281250
   "001111000110010000", -- Line 1   Column 1046   Coefficient 60.39062500
   "001111000110011001", -- Line 1   Column 1047   Coefficient 60.39941406
   "001111000110100001", -- Line 1   Column 1048   Coefficient 60.40722656
   "001111000110101001", -- Line 1   Column 1049   Coefficient 60.41503906
   "001111000110110010", -- Line 1   Column 1050   Coefficient 60.42382813
   "001111000110111010", -- Line 1   Column 1051   Coefficient 60.43164063
   "001111000111000011", -- Line 1   Column 1052   Coefficient 60.44042969
   "001111000111001011", -- Line 1   Column 1053   Coefficient 60.44824219
   "001111000111010100", -- Line 1   Column 1054   Coefficient 60.45703125
   "001111000111011100", -- Line 1   Column 1055   Coefficient 60.46484375
   "001111000111100101", -- Line 1   Column 1056   Coefficient 60.47363281
   "001111000111101101", -- Line 1   Column 1057   Coefficient 60.48144531
   "001111000111110101", -- Line 1   Column 1058   Coefficient 60.48925781
   "001111000111111110", -- Line 1   Column 1059   Coefficient 60.49804688
   "001111001000000110", -- Line 1   Column 1060   Coefficient 60.50585938
   "001111001000001111", -- Line 1   Column 1061   Coefficient 60.51464844
   "001111001000010111", -- Line 1   Column 1062   Coefficient 60.52246094
   "001111001000011111", -- Line 1   Column 1063   Coefficient 60.53027344
   "001111001000101000", -- Line 1   Column 1064   Coefficient 60.53906250
   "001111001000110000", -- Line 1   Column 1065   Coefficient 60.54687500
   "001111001000111000", -- Line 1   Column 1066   Coefficient 60.55468750
   "001111001001000001", -- Line 1   Column 1067   Coefficient 60.56347656
   "001111001001001001", -- Line 1   Column 1068   Coefficient 60.57128906
   "001111001001010001", -- Line 1   Column 1069   Coefficient 60.57910156
   "001111001001011010", -- Line 1   Column 1070   Coefficient 60.58789063
   "001111001001100010", -- Line 1   Column 1071   Coefficient 60.59570313
   "001111001001101010", -- Line 1   Column 1072   Coefficient 60.60351563
   "001111001001110011", -- Line 1   Column 1073   Coefficient 60.61230469
   "001111001001111011", -- Line 1   Column 1074   Coefficient 60.62011719
   "001111001010000011", -- Line 1   Column 1075   Coefficient 60.62792969
   "001111001010001100", -- Line 1   Column 1076   Coefficient 60.63671875
   "001111001010010100", -- Line 1   Column 1077   Coefficient 60.64453125
   "001111001010011100", -- Line 1   Column 1078   Coefficient 60.65234375
   "001111001010100100", -- Line 1   Column 1079   Coefficient 60.66015625
   "001111001010101101", -- Line 1   Column 1080   Coefficient 60.66894531
   "001111001010110101", -- Line 1   Column 1081   Coefficient 60.67675781
   "001111001010111101", -- Line 1   Column 1082   Coefficient 60.68457031
   "001111001011000101", -- Line 1   Column 1083   Coefficient 60.69238281
   "001111001011001101", -- Line 1   Column 1084   Coefficient 60.70019531
   "001111001011010110", -- Line 1   Column 1085   Coefficient 60.70898438
   "001111001011011110", -- Line 1   Column 1086   Coefficient 60.71679688
   "001111001011100110", -- Line 1   Column 1087   Coefficient 60.72460938
   "001111001011101110", -- Line 1   Column 1088   Coefficient 60.73242188
   "001111001011110110", -- Line 1   Column 1089   Coefficient 60.74023438
   "001111001011111110", -- Line 1   Column 1090   Coefficient 60.74804688
   "001111001100000111", -- Line 1   Column 1091   Coefficient 60.75683594
   "001111001100001111", -- Line 1   Column 1092   Coefficient 60.76464844
   "001111001100010111", -- Line 1   Column 1093   Coefficient 60.77246094
   "001111001100011111", -- Line 1   Column 1094   Coefficient 60.78027344
   "001111001100100111", -- Line 1   Column 1095   Coefficient 60.78808594
   "001111001100101111", -- Line 1   Column 1096   Coefficient 60.79589844
   "001111001100110111", -- Line 1   Column 1097   Coefficient 60.80371094
   "001111001101000000", -- Line 1   Column 1098   Coefficient 60.81250000
   "001111001101001000", -- Line 1   Column 1099   Coefficient 60.82031250
   "001111001101010000", -- Line 1   Column 1100   Coefficient 60.82812500
   "001111001101011000", -- Line 1   Column 1101   Coefficient 60.83593750
   "001111001101100000", -- Line 1   Column 1102   Coefficient 60.84375000
   "001111001101101000", -- Line 1   Column 1103   Coefficient 60.85156250
   "001111001101110000", -- Line 1   Column 1104   Coefficient 60.85937500
   "001111001101111000", -- Line 1   Column 1105   Coefficient 60.86718750
   "001111001110000000", -- Line 1   Column 1106   Coefficient 60.87500000
   "001111001110001000", -- Line 1   Column 1107   Coefficient 60.88281250
   "001111001110010000", -- Line 1   Column 1108   Coefficient 60.89062500
   "001111001110011000", -- Line 1   Column 1109   Coefficient 60.89843750
   "001111001110100000", -- Line 1   Column 1110   Coefficient 60.90625000
   "001111001110101000", -- Line 1   Column 1111   Coefficient 60.91406250
   "001111001110110000", -- Line 1   Column 1112   Coefficient 60.92187500
   "001111001110111000", -- Line 1   Column 1113   Coefficient 60.92968750
   "001111001111000000", -- Line 1   Column 1114   Coefficient 60.93750000
   "001111001111001000", -- Line 1   Column 1115   Coefficient 60.94531250
   "001111001111010000", -- Line 1   Column 1116   Coefficient 60.95312500
   "001111001111011000", -- Line 1   Column 1117   Coefficient 60.96093750
   "001111001111100000", -- Line 1   Column 1118   Coefficient 60.96875000
   "001111001111101000", -- Line 1   Column 1119   Coefficient 60.97656250
   "001111001111110000", -- Line 1   Column 1120   Coefficient 60.98437500
   "001111001111111000", -- Line 1   Column 1121   Coefficient 60.99218750
   "001111010000000000", -- Line 1   Column 1122   Coefficient 61.00000000
   "001111010000001000", -- Line 1   Column 1123   Coefficient 61.00781250
   "001111010000010000", -- Line 1   Column 1124   Coefficient 61.01562500
   "001111010000011000", -- Line 1   Column 1125   Coefficient 61.02343750
   "001111010000100000", -- Line 1   Column 1126   Coefficient 61.03125000
   "001111010000100111", -- Line 1   Column 1127   Coefficient 61.03808594
   "001111010000101111", -- Line 1   Column 1128   Coefficient 61.04589844
   "001111010000110111", -- Line 1   Column 1129   Coefficient 61.05371094
   "001111010000111111", -- Line 1   Column 1130   Coefficient 61.06152344
   "001111010001000111", -- Line 1   Column 1131   Coefficient 61.06933594
   "001111010001001111", -- Line 1   Column 1132   Coefficient 61.07714844
   "001111010001010111", -- Line 1   Column 1133   Coefficient 61.08496094
   "001111010001011110", -- Line 1   Column 1134   Coefficient 61.09179688
   "001111010001100110", -- Line 1   Column 1135   Coefficient 61.09960938
   "001111010001101110", -- Line 1   Column 1136   Coefficient 61.10742188
   "001111010001110110", -- Line 1   Column 1137   Coefficient 61.11523438
   "001111010001111110", -- Line 1   Column 1138   Coefficient 61.12304688
   "001111010010000110", -- Line 1   Column 1139   Coefficient 61.13085938
   "001111010010001101", -- Line 1   Column 1140   Coefficient 61.13769531
   "001111010010010101", -- Line 1   Column 1141   Coefficient 61.14550781
   "001111010010011101", -- Line 1   Column 1142   Coefficient 61.15332031
   "001111010010100101", -- Line 1   Column 1143   Coefficient 61.16113281
   "001111010010101101", -- Line 1   Column 1144   Coefficient 61.16894531
   "001111010010110100", -- Line 1   Column 1145   Coefficient 61.17578125
   "001111010010111100", -- Line 1   Column 1146   Coefficient 61.18359375
   "001111010011000100", -- Line 1   Column 1147   Coefficient 61.19140625
   "001111010011001100", -- Line 1   Column 1148   Coefficient 61.19921875
   "001111010011010011", -- Line 1   Column 1149   Coefficient 61.20605469
   "001111010011011011", -- Line 1   Column 1150   Coefficient 61.21386719
   "001111010011100011", -- Line 1   Column 1151   Coefficient 61.22167969
   "001111010011101011", -- Line 1   Column 1152   Coefficient 61.22949219
   "001111010011110010", -- Line 1   Column 1153   Coefficient 61.23632813
   "001111010011111010", -- Line 1   Column 1154   Coefficient 61.24414063
   "001111010100000010", -- Line 1   Column 1155   Coefficient 61.25195313
   "001111010100001001", -- Line 1   Column 1156   Coefficient 61.25878906
   "001111010100010001", -- Line 1   Column 1157   Coefficient 61.26660156
   "001111010100011001", -- Line 1   Column 1158   Coefficient 61.27441406
   "001111010100100000", -- Line 1   Column 1159   Coefficient 61.28125000
   "001111010100101000", -- Line 1   Column 1160   Coefficient 61.28906250
   "001111010100110000", -- Line 1   Column 1161   Coefficient 61.29687500
   "001111010100110111", -- Line 1   Column 1162   Coefficient 61.30371094
   "001111010100111111", -- Line 1   Column 1163   Coefficient 61.31152344
   "001111010101000111", -- Line 1   Column 1164   Coefficient 61.31933594
   "001111010101001110", -- Line 1   Column 1165   Coefficient 61.32617188
   "001111010101010110", -- Line 1   Column 1166   Coefficient 61.33398438
   "001111010101011110", -- Line 1   Column 1167   Coefficient 61.34179688
   "001111010101100101", -- Line 1   Column 1168   Coefficient 61.34863281
   "001111010101101101", -- Line 1   Column 1169   Coefficient 61.35644531
   "001111010101110100", -- Line 1   Column 1170   Coefficient 61.36328125
   "001111010101111100", -- Line 1   Column 1171   Coefficient 61.37109375
   "001111010110000100", -- Line 1   Column 1172   Coefficient 61.37890625
   "001111010110001011", -- Line 1   Column 1173   Coefficient 61.38574219
   "001111010110010011", -- Line 1   Column 1174   Coefficient 61.39355469
   "001111010110011010", -- Line 1   Column 1175   Coefficient 61.40039063
   "001111010110100010", -- Line 1   Column 1176   Coefficient 61.40820313
   "001111010110101010", -- Line 1   Column 1177   Coefficient 61.41601563
   "001111010110110001", -- Line 1   Column 1178   Coefficient 61.42285156
   "001111010110111001", -- Line 1   Column 1179   Coefficient 61.43066406
   "001111010111000000", -- Line 1   Column 1180   Coefficient 61.43750000
   "001111010111001000", -- Line 1   Column 1181   Coefficient 61.44531250
   "001111010111001111", -- Line 1   Column 1182   Coefficient 61.45214844
   "001111010111010111", -- Line 1   Column 1183   Coefficient 61.45996094
   "001111010111011110", -- Line 1   Column 1184   Coefficient 61.46679688
   "001111010111100110", -- Line 1   Column 1185   Coefficient 61.47460938
   "001111010111101101", -- Line 1   Column 1186   Coefficient 61.48144531
   "001111010111110101", -- Line 1   Column 1187   Coefficient 61.48925781
   "001111010111111100", -- Line 1   Column 1188   Coefficient 61.49609375
   "001111011000000100", -- Line 1   Column 1189   Coefficient 61.50390625
   "001111011000001011", -- Line 1   Column 1190   Coefficient 61.51074219
   "001111011000010011", -- Line 1   Column 1191   Coefficient 61.51855469
   "001111011000011010", -- Line 1   Column 1192   Coefficient 61.52539063
   "001111011000100010", -- Line 1   Column 1193   Coefficient 61.53320313
   "001111011000101001", -- Line 1   Column 1194   Coefficient 61.54003906
   "001111011000110000", -- Line 1   Column 1195   Coefficient 61.54687500
   "001111011000111000", -- Line 1   Column 1196   Coefficient 61.55468750
   "001111011000111111", -- Line 1   Column 1197   Coefficient 61.56152344
   "001111011001000111", -- Line 1   Column 1198   Coefficient 61.56933594
   "001111011001001110", -- Line 1   Column 1199   Coefficient 61.57617188
   "001111011001010110", -- Line 1   Column 1200   Coefficient 61.58398438
   "001111011001011101", -- Line 1   Column 1201   Coefficient 61.59082031
   "001111011001100100", -- Line 1   Column 1202   Coefficient 61.59765625
   "001111011001101100", -- Line 1   Column 1203   Coefficient 61.60546875
   "001111011001110011", -- Line 1   Column 1204   Coefficient 61.61230469
   "001111011001111011", -- Line 1   Column 1205   Coefficient 61.62011719
   "001111011010000010", -- Line 1   Column 1206   Coefficient 61.62695313
   "001111011010001001", -- Line 1   Column 1207   Coefficient 61.63378906
   "001111011010010001", -- Line 1   Column 1208   Coefficient 61.64160156
   "001111011010011000", -- Line 1   Column 1209   Coefficient 61.64843750
   "001111011010011111", -- Line 1   Column 1210   Coefficient 61.65527344
   "001111011010100111", -- Line 1   Column 1211   Coefficient 61.66308594
   "001111011010101110", -- Line 1   Column 1212   Coefficient 61.66992188
   "001111011010110101", -- Line 1   Column 1213   Coefficient 61.67675781
   "001111011010111101", -- Line 1   Column 1214   Coefficient 61.68457031
   "001111011011000100", -- Line 1   Column 1215   Coefficient 61.69140625
   "001111011011001011", -- Line 1   Column 1216   Coefficient 61.69824219
   "001111011011010011", -- Line 1   Column 1217   Coefficient 61.70605469
   "001111011011011010", -- Line 1   Column 1218   Coefficient 61.71289063
   "001111011011100001", -- Line 1   Column 1219   Coefficient 61.71972656
   "001111011011101001", -- Line 1   Column 1220   Coefficient 61.72753906
   "001111011011110000", -- Line 1   Column 1221   Coefficient 61.73437500
   "001111011011110111", -- Line 1   Column 1222   Coefficient 61.74121094
   "001111011011111110", -- Line 1   Column 1223   Coefficient 61.74804688
   "001111011100000110", -- Line 1   Column 1224   Coefficient 61.75585938
   "001111011100001101", -- Line 1   Column 1225   Coefficient 61.76269531
   "001111011100010100", -- Line 1   Column 1226   Coefficient 61.76953125
   "001111011100011100", -- Line 1   Column 1227   Coefficient 61.77734375
   "001111011100100011", -- Line 1   Column 1228   Coefficient 61.78417969
   "001111011100101010", -- Line 1   Column 1229   Coefficient 61.79101563
   "001111011100110001", -- Line 1   Column 1230   Coefficient 61.79785156
   "001111011100111000", -- Line 1   Column 1231   Coefficient 61.80468750
   "001111011101000000", -- Line 1   Column 1232   Coefficient 61.81250000
   "001111011101000111", -- Line 1   Column 1233   Coefficient 61.81933594
   "001111011101001110", -- Line 1   Column 1234   Coefficient 61.82617188
   "001111011101010101", -- Line 1   Column 1235   Coefficient 61.83300781
   "001111011101011101", -- Line 1   Column 1236   Coefficient 61.84082031
   "001111011101100100", -- Line 1   Column 1237   Coefficient 61.84765625
   "001111011101101011", -- Line 1   Column 1238   Coefficient 61.85449219
   "001111011101110010", -- Line 1   Column 1239   Coefficient 61.86132813
   "001111011101111001", -- Line 1   Column 1240   Coefficient 61.86816406
   "001111011110000000", -- Line 1   Column 1241   Coefficient 61.87500000
   "001111011110001000", -- Line 1   Column 1242   Coefficient 61.88281250
   "001111011110001111", -- Line 1   Column 1243   Coefficient 61.88964844
   "001111011110010110", -- Line 1   Column 1244   Coefficient 61.89648438
   "001111011110011101", -- Line 1   Column 1245   Coefficient 61.90332031
   "001111011110100100", -- Line 1   Column 1246   Coefficient 61.91015625
   "001111011110101011", -- Line 1   Column 1247   Coefficient 61.91699219
   "001111011110110010", -- Line 1   Column 1248   Coefficient 61.92382813
   "001111011110111010", -- Line 1   Column 1249   Coefficient 61.93164063
   "001111011111000001", -- Line 1   Column 1250   Coefficient 61.93847656
   "001111011111001000", -- Line 1   Column 1251   Coefficient 61.94531250
   "001111011111001111", -- Line 1   Column 1252   Coefficient 61.95214844
   "001111011111010110", -- Line 1   Column 1253   Coefficient 61.95898438
   "001111011111011101", -- Line 1   Column 1254   Coefficient 61.96582031
   "001111011111100100", -- Line 1   Column 1255   Coefficient 61.97265625
   "001111011111101011", -- Line 1   Column 1256   Coefficient 61.97949219
   "001111011111110010", -- Line 1   Column 1257   Coefficient 61.98632813
   "001111011111111001", -- Line 1   Column 1258   Coefficient 61.99316406
   "001111100000000001", -- Line 1   Column 1259   Coefficient 62.00097656
   "001111100000001000", -- Line 1   Column 1260   Coefficient 62.00781250
   "001111100000001111", -- Line 1   Column 1261   Coefficient 62.01464844
   "001111100000010110", -- Line 1   Column 1262   Coefficient 62.02148438
   "001111100000011101", -- Line 1   Column 1263   Coefficient 62.02832031
   "001111100000100100", -- Line 1   Column 1264   Coefficient 62.03515625
   "001111100000101011", -- Line 1   Column 1265   Coefficient 62.04199219
   "001111100000110010", -- Line 1   Column 1266   Coefficient 62.04882813
   "001111100000111001", -- Line 1   Column 1267   Coefficient 62.05566406
   "001111100001000000", -- Line 1   Column 1268   Coefficient 62.06250000
   "001111100001000111", -- Line 1   Column 1269   Coefficient 62.06933594
   "001111100001001110", -- Line 1   Column 1270   Coefficient 62.07617188
   "001111100001010101", -- Line 1   Column 1271   Coefficient 62.08300781
   "001111100001011100", -- Line 1   Column 1272   Coefficient 62.08984375
   "001111100001100011", -- Line 1   Column 1273   Coefficient 62.09667969
   "001111100001101010", -- Line 1   Column 1274   Coefficient 62.10351563
   "001111100001110001", -- Line 1   Column 1275   Coefficient 62.11035156
   "001111100001111000", -- Line 1   Column 1276   Coefficient 62.11718750
   "001111100001111111", -- Line 1   Column 1277   Coefficient 62.12402344
   "001111100010000110", -- Line 1   Column 1278   Coefficient 62.13085938
   "001111100010001101", -- Line 1   Column 1279   Coefficient 62.13769531
   "001111100010010100", -- Line 1   Column 1280   Coefficient 62.14453125
   "001111100010011011", -- Line 1   Column 1281   Coefficient 62.15136719
   "001111100010100010", -- Line 1   Column 1282   Coefficient 62.15820313
   "001111100010101000", -- Line 1   Column 1283   Coefficient 62.16406250
   "001111100010101111", -- Line 1   Column 1284   Coefficient 62.17089844
   "001111100010110110", -- Line 1   Column 1285   Coefficient 62.17773438
   "001111100010111101", -- Line 1   Column 1286   Coefficient 62.18457031
   "001111100011000100", -- Line 1   Column 1287   Coefficient 62.19140625
   "001111100011001011", -- Line 1   Column 1288   Coefficient 62.19824219
   "001111100011010010", -- Line 1   Column 1289   Coefficient 62.20507813
   "001111100011011001", -- Line 1   Column 1290   Coefficient 62.21191406
   "001111100011100000", -- Line 1   Column 1291   Coefficient 62.21875000
   "001111100011100111", -- Line 1   Column 1292   Coefficient 62.22558594
   "001111100011101110", -- Line 1   Column 1293   Coefficient 62.23242188
   "001111100011110100", -- Line 1   Column 1294   Coefficient 62.23828125
   "001111100011111011", -- Line 1   Column 1295   Coefficient 62.24511719
   "001111100100000010", -- Line 1   Column 1296   Coefficient 62.25195313
   "001111100100001001", -- Line 1   Column 1297   Coefficient 62.25878906
   "001111100100010000", -- Line 1   Column 1298   Coefficient 62.26562500
   "001111100100010111", -- Line 1   Column 1299   Coefficient 62.27246094
   "001111100100011110", -- Line 1   Column 1300   Coefficient 62.27929688
   "001111100100100100", -- Line 1   Column 1301   Coefficient 62.28515625
   "001111100100101011", -- Line 1   Column 1302   Coefficient 62.29199219
   "001111100100110010", -- Line 1   Column 1303   Coefficient 62.29882813
   "001111100100111001", -- Line 1   Column 1304   Coefficient 62.30566406
   "001111100101000000", -- Line 1   Column 1305   Coefficient 62.31250000
   "001111100101000111", -- Line 1   Column 1306   Coefficient 62.31933594
   "001111100101001101", -- Line 1   Column 1307   Coefficient 62.32519531
   "001111100101010100", -- Line 1   Column 1308   Coefficient 62.33203125
   "001111100101011011", -- Line 1   Column 1309   Coefficient 62.33886719
   "001111100101100010", -- Line 1   Column 1310   Coefficient 62.34570313
   "001111100101101001", -- Line 1   Column 1311   Coefficient 62.35253906
   "001111100101101111", -- Line 1   Column 1312   Coefficient 62.35839844
   "001111100101110110", -- Line 1   Column 1313   Coefficient 62.36523438
   "001111100101111101", -- Line 1   Column 1314   Coefficient 62.37207031
   "001111100110000100", -- Line 1   Column 1315   Coefficient 62.37890625
   "001111100110001010", -- Line 1   Column 1316   Coefficient 62.38476563
   "001111100110010001", -- Line 1   Column 1317   Coefficient 62.39160156
   "001111100110011000", -- Line 1   Column 1318   Coefficient 62.39843750
   "001111100110011111", -- Line 1   Column 1319   Coefficient 62.40527344
   "001111100110100101", -- Line 1   Column 1320   Coefficient 62.41113281
   "001111100110101100", -- Line 1   Column 1321   Coefficient 62.41796875
   "001111100110110011", -- Line 1   Column 1322   Coefficient 62.42480469
   "001111100110111010", -- Line 1   Column 1323   Coefficient 62.43164063
   "001111100111000000", -- Line 1   Column 1324   Coefficient 62.43750000
   "001111100111000111", -- Line 1   Column 1325   Coefficient 62.44433594
   "001111100111001110", -- Line 1   Column 1326   Coefficient 62.45117188
   "001111100111010100", -- Line 1   Column 1327   Coefficient 62.45703125
   "001111100111011011", -- Line 1   Column 1328   Coefficient 62.46386719
   "001111100111100010", -- Line 1   Column 1329   Coefficient 62.47070313
   "001111100111101000", -- Line 1   Column 1330   Coefficient 62.47656250
   "001111100111101111", -- Line 1   Column 1331   Coefficient 62.48339844
   "001111100111110110", -- Line 1   Column 1332   Coefficient 62.49023438
   "001111100111111101", -- Line 1   Column 1333   Coefficient 62.49707031
   "001111101000000011", -- Line 1   Column 1334   Coefficient 62.50292969
   "001111101000001010", -- Line 1   Column 1335   Coefficient 62.50976563
   "001111101000010001", -- Line 1   Column 1336   Coefficient 62.51660156
   "001111101000010111", -- Line 1   Column 1337   Coefficient 62.52246094
   "001111101000011110", -- Line 1   Column 1338   Coefficient 62.52929688
   "001111101000100100", -- Line 1   Column 1339   Coefficient 62.53515625
   "001111101000101011", -- Line 1   Column 1340   Coefficient 62.54199219
   "001111101000110010", -- Line 1   Column 1341   Coefficient 62.54882813
   "001111101000111000", -- Line 1   Column 1342   Coefficient 62.55468750
   "001111101000111111", -- Line 1   Column 1343   Coefficient 62.56152344
   "001111101001000110", -- Line 1   Column 1344   Coefficient 62.56835938
   "001111101001001100", -- Line 1   Column 1345   Coefficient 62.57421875
   "001111101001010011", -- Line 1   Column 1346   Coefficient 62.58105469
   "001111101001011001", -- Line 1   Column 1347   Coefficient 62.58691406
   "001111101001100000", -- Line 1   Column 1348   Coefficient 62.59375000
   "001111101001100111", -- Line 1   Column 1349   Coefficient 62.60058594
   "001111101001101101", -- Line 1   Column 1350   Coefficient 62.60644531
   "001111101001110100", -- Line 1   Column 1351   Coefficient 62.61328125
   "001111101001111010", -- Line 1   Column 1352   Coefficient 62.61914063
   "001111101010000001", -- Line 1   Column 1353   Coefficient 62.62597656
   "001111101010001000", -- Line 1   Column 1354   Coefficient 62.63281250
   "001111101010001110", -- Line 1   Column 1355   Coefficient 62.63867188
   "001111101010010101", -- Line 1   Column 1356   Coefficient 62.64550781
   "001111101010011011", -- Line 1   Column 1357   Coefficient 62.65136719
   "001111101010100010", -- Line 1   Column 1358   Coefficient 62.65820313
   "001111101010101000", -- Line 1   Column 1359   Coefficient 62.66406250
   "001111101010101111", -- Line 1   Column 1360   Coefficient 62.67089844
   "001111101010110101", -- Line 1   Column 1361   Coefficient 62.67675781
   "001111101010111100", -- Line 1   Column 1362   Coefficient 62.68359375
   "001111101011000010", -- Line 1   Column 1363   Coefficient 62.68945313
   "001111101011001001", -- Line 1   Column 1364   Coefficient 62.69628906
   "001111101011010000", -- Line 1   Column 1365   Coefficient 62.70312500
   "001111101011010110", -- Line 1   Column 1366   Coefficient 62.70898438
   "001111101011011101", -- Line 1   Column 1367   Coefficient 62.71582031
   "001111101011100011", -- Line 1   Column 1368   Coefficient 62.72167969
   "001111101011101010", -- Line 1   Column 1369   Coefficient 62.72851563
   "001111101011110000", -- Line 1   Column 1370   Coefficient 62.73437500
   "001111101011110111", -- Line 1   Column 1371   Coefficient 62.74121094
   "001111101011111101", -- Line 1   Column 1372   Coefficient 62.74707031
   "001111101100000011", -- Line 1   Column 1373   Coefficient 62.75292969
   "001111101100001010", -- Line 1   Column 1374   Coefficient 62.75976563
   "001111101100010000", -- Line 1   Column 1375   Coefficient 62.76562500
   "001111101100010111", -- Line 1   Column 1376   Coefficient 62.77246094
   "001111101100011101", -- Line 1   Column 1377   Coefficient 62.77832031
   "001111101100100100", -- Line 1   Column 1378   Coefficient 62.78515625
   "001111101100101010", -- Line 1   Column 1379   Coefficient 62.79101563
   "001111101100110001", -- Line 1   Column 1380   Coefficient 62.79785156
   "001111101100110111", -- Line 1   Column 1381   Coefficient 62.80371094
   "001111101100111110", -- Line 1   Column 1382   Coefficient 62.81054688
   "001111101101000100", -- Line 1   Column 1383   Coefficient 62.81640625
   "001111101101001010", -- Line 1   Column 1384   Coefficient 62.82226563
   "001111101101010001", -- Line 1   Column 1385   Coefficient 62.82910156
   "001111101101010111", -- Line 1   Column 1386   Coefficient 62.83496094
   "001111101101011110", -- Line 1   Column 1387   Coefficient 62.84179688
   "001111101101100100", -- Line 1   Column 1388   Coefficient 62.84765625
   "001111101101101011", -- Line 1   Column 1389   Coefficient 62.85449219
   "001111101101110001", -- Line 1   Column 1390   Coefficient 62.86035156
   "001111101101110111", -- Line 1   Column 1391   Coefficient 62.86621094
   "001111101101111110", -- Line 1   Column 1392   Coefficient 62.87304688
   "001111101110000100", -- Line 1   Column 1393   Coefficient 62.87890625
   "001111101110001011", -- Line 1   Column 1394   Coefficient 62.88574219
   "001111101110010001", -- Line 1   Column 1395   Coefficient 62.89160156
   "001111101110010111", -- Line 1   Column 1396   Coefficient 62.89746094
   "001111101110011110", -- Line 1   Column 1397   Coefficient 62.90429688
   "001111101110100100", -- Line 1   Column 1398   Coefficient 62.91015625
   "001111101110101010", -- Line 1   Column 1399   Coefficient 62.91601563
   "001111101110110001", -- Line 1   Column 1400   Coefficient 62.92285156
   "001111101110110111", -- Line 1   Column 1401   Coefficient 62.92871094
   "001111101110111101", -- Line 1   Column 1402   Coefficient 62.93457031
   "001111101111000100", -- Line 1   Column 1403   Coefficient 62.94140625
   "001111101111001010", -- Line 1   Column 1404   Coefficient 62.94726563
   "001111101111010000", -- Line 1   Column 1405   Coefficient 62.95312500
   "001111101111010111", -- Line 1   Column 1406   Coefficient 62.95996094
   "001111101111011101", -- Line 1   Column 1407   Coefficient 62.96582031
   "001111101111100011", -- Line 1   Column 1408   Coefficient 62.97167969
   "001111101111101010", -- Line 1   Column 1409   Coefficient 62.97851563
   "001111101111110000", -- Line 1   Column 1410   Coefficient 62.98437500
   "001111101111110110", -- Line 1   Column 1411   Coefficient 62.99023438
   "001111101111111101", -- Line 1   Column 1412   Coefficient 62.99707031
   "001111110000000011", -- Line 1   Column 1413   Coefficient 63.00292969
   "001111110000001001", -- Line 1   Column 1414   Coefficient 63.00878906
   "001111110000001111", -- Line 1   Column 1415   Coefficient 63.01464844
   "001111110000010110", -- Line 1   Column 1416   Coefficient 63.02148438
   "001111110000011100", -- Line 1   Column 1417   Coefficient 63.02734375
   "001111110000100010", -- Line 1   Column 1418   Coefficient 63.03320313
   "001111110000101001", -- Line 1   Column 1419   Coefficient 63.04003906
   "001111110000101111", -- Line 1   Column 1420   Coefficient 63.04589844
   "001111110000110101", -- Line 1   Column 1421   Coefficient 63.05175781
   "001111110000111011", -- Line 1   Column 1422   Coefficient 63.05761719
   "001111110001000010", -- Line 1   Column 1423   Coefficient 63.06445313
   "001111110001001000", -- Line 1   Column 1424   Coefficient 63.07031250
   "001111110001001110", -- Line 1   Column 1425   Coefficient 63.07617188
   "001111110001010100", -- Line 1   Column 1426   Coefficient 63.08203125
   "001111110001011011", -- Line 1   Column 1427   Coefficient 63.08886719
   "001111110001100001", -- Line 1   Column 1428   Coefficient 63.09472656
   "001111110001100111", -- Line 1   Column 1429   Coefficient 63.10058594
   "001111110001101101", -- Line 1   Column 1430   Coefficient 63.10644531
   "001111110001110011", -- Line 1   Column 1431   Coefficient 63.11230469
   "001111110001111010", -- Line 1   Column 1432   Coefficient 63.11914063
   "001111110010000000", -- Line 1   Column 1433   Coefficient 63.12500000
   "001111110010000110", -- Line 1   Column 1434   Coefficient 63.13085938
   "001111110010001100", -- Line 1   Column 1435   Coefficient 63.13671875
   "001111110010010011", -- Line 1   Column 1436   Coefficient 63.14355469
   "001111110010011001", -- Line 1   Column 1437   Coefficient 63.14941406
   "001111110010011111", -- Line 1   Column 1438   Coefficient 63.15527344
   "001111110010100101", -- Line 1   Column 1439   Coefficient 63.16113281
   "001111110010101011", -- Line 1   Column 1440   Coefficient 63.16699219
   "001111110010110001", -- Line 1   Column 1441   Coefficient 63.17285156
   "001111110010111000", -- Line 1   Column 1442   Coefficient 63.17968750
   "001111110010111110", -- Line 1   Column 1443   Coefficient 63.18554688
   "001111110011000100", -- Line 1   Column 1444   Coefficient 63.19140625
   "001111110011001010", -- Line 1   Column 1445   Coefficient 63.19726563
   "001111110011010000", -- Line 1   Column 1446   Coefficient 63.20312500
   "001111110011010110", -- Line 1   Column 1447   Coefficient 63.20898438
   "001111110011011101", -- Line 1   Column 1448   Coefficient 63.21582031
   "001111110011100011", -- Line 1   Column 1449   Coefficient 63.22167969
   "001111110011101001", -- Line 1   Column 1450   Coefficient 63.22753906
   "001111110011101111", -- Line 1   Column 1451   Coefficient 63.23339844
   "001111110011110101", -- Line 1   Column 1452   Coefficient 63.23925781
   "001111110011111011", -- Line 1   Column 1453   Coefficient 63.24511719
   "001111110100000001", -- Line 1   Column 1454   Coefficient 63.25097656
   "001111110100000111", -- Line 1   Column 1455   Coefficient 63.25683594
   "001111110100001110", -- Line 1   Column 1456   Coefficient 63.26367188
   "001111110100010100", -- Line 1   Column 1457   Coefficient 63.26953125
   "001111110100011010", -- Line 1   Column 1458   Coefficient 63.27539063
   "001111110100100000", -- Line 1   Column 1459   Coefficient 63.28125000
   "001111110100100110", -- Line 1   Column 1460   Coefficient 63.28710938
   "001111110100101100", -- Line 1   Column 1461   Coefficient 63.29296875
   "001111110100110010", -- Line 1   Column 1462   Coefficient 63.29882813
   "001111110100111000", -- Line 1   Column 1463   Coefficient 63.30468750
   "001111110100111110", -- Line 1   Column 1464   Coefficient 63.31054688
   "001111110101000100", -- Line 1   Column 1465   Coefficient 63.31640625
   "001111110101001010", -- Line 1   Column 1466   Coefficient 63.32226563
   "001111110101010000", -- Line 1   Column 1467   Coefficient 63.32812500
   "001111110101010111", -- Line 1   Column 1468   Coefficient 63.33496094
   "001111110101011101", -- Line 1   Column 1469   Coefficient 63.34082031
   "001111110101100011", -- Line 1   Column 1470   Coefficient 63.34667969
   "001111110101101001", -- Line 1   Column 1471   Coefficient 63.35253906
   "001111110101101111", -- Line 1   Column 1472   Coefficient 63.35839844
   "001111110101110101", -- Line 1   Column 1473   Coefficient 63.36425781
   "001111110101111011", -- Line 1   Column 1474   Coefficient 63.37011719
   "001111110110000001", -- Line 1   Column 1475   Coefficient 63.37597656
   "001111110110000111", -- Line 1   Column 1476   Coefficient 63.38183594
   "001111110110001101", -- Line 1   Column 1477   Coefficient 63.38769531
   "001111110110010011", -- Line 1   Column 1478   Coefficient 63.39355469
   "001111110110011001", -- Line 1   Column 1479   Coefficient 63.39941406
   "001111110110011111", -- Line 1   Column 1480   Coefficient 63.40527344
   "001111110110100101", -- Line 1   Column 1481   Coefficient 63.41113281
   "001111110110101011", -- Line 1   Column 1482   Coefficient 63.41699219
   "001111110110110001", -- Line 1   Column 1483   Coefficient 63.42285156
   "001111110110110111", -- Line 1   Column 1484   Coefficient 63.42871094
   "001111110110111101", -- Line 1   Column 1485   Coefficient 63.43457031
   "001111110111000011", -- Line 1   Column 1486   Coefficient 63.44042969
   "001111110111001001", -- Line 1   Column 1487   Coefficient 63.44628906
   "001111110111001111", -- Line 1   Column 1488   Coefficient 63.45214844
   "001111110111010101", -- Line 1   Column 1489   Coefficient 63.45800781
   "001111110111011011", -- Line 1   Column 1490   Coefficient 63.46386719
   "001111110111100001", -- Line 1   Column 1491   Coefficient 63.46972656
   "001111110111100111", -- Line 1   Column 1492   Coefficient 63.47558594
   "001111110111101101", -- Line 1   Column 1493   Coefficient 63.48144531
   "001111110111110011", -- Line 1   Column 1494   Coefficient 63.48730469
   "001111110111111001", -- Line 1   Column 1495   Coefficient 63.49316406
   "001111110111111111", -- Line 1   Column 1496   Coefficient 63.49902344
   "001111111000000101", -- Line 1   Column 1497   Coefficient 63.50488281
   "001111111000001010", -- Line 1   Column 1498   Coefficient 63.50976563
   "001111111000010000", -- Line 1   Column 1499   Coefficient 63.51562500
   "001111111000010110", -- Line 1   Column 1500   Coefficient 63.52148438
   "001111111000011100", -- Line 1   Column 1501   Coefficient 63.52734375
   "001111111000100010", -- Line 1   Column 1502   Coefficient 63.53320313
   "001111111000101000", -- Line 1   Column 1503   Coefficient 63.53906250
   "001111111000101110", -- Line 1   Column 1504   Coefficient 63.54492188
   "001111111000110100", -- Line 1   Column 1505   Coefficient 63.55078125
   "001111111000111010", -- Line 1   Column 1506   Coefficient 63.55664063
   "001111111001000000", -- Line 1   Column 1507   Coefficient 63.56250000
   "001111111001000110", -- Line 1   Column 1508   Coefficient 63.56835938
   "001111111001001100", -- Line 1   Column 1509   Coefficient 63.57421875
   "001111111001010001", -- Line 1   Column 1510   Coefficient 63.57910156
   "001111111001010111", -- Line 1   Column 1511   Coefficient 63.58496094
   "001111111001011101", -- Line 1   Column 1512   Coefficient 63.59082031
   "001111111001100011", -- Line 1   Column 1513   Coefficient 63.59667969
   "001111111001101001", -- Line 1   Column 1514   Coefficient 63.60253906
   "001111111001101111", -- Line 1   Column 1515   Coefficient 63.60839844
   "001111111001110101", -- Line 1   Column 1516   Coefficient 63.61425781
   "001111111001111011", -- Line 1   Column 1517   Coefficient 63.62011719
   "001111111010000000", -- Line 1   Column 1518   Coefficient 63.62500000
   "001111111010000110", -- Line 1   Column 1519   Coefficient 63.63085938
   "001111111010001100", -- Line 1   Column 1520   Coefficient 63.63671875
   "001111111010010010", -- Line 1   Column 1521   Coefficient 63.64257813
   "001111111010011000", -- Line 1   Column 1522   Coefficient 63.64843750
   "001111111010011110", -- Line 1   Column 1523   Coefficient 63.65429688
   "001111111010100100", -- Line 1   Column 1524   Coefficient 63.66015625
   "001111111010101001", -- Line 1   Column 1525   Coefficient 63.66503906
   "001111111010101111", -- Line 1   Column 1526   Coefficient 63.67089844
   "001111111010110101", -- Line 1   Column 1527   Coefficient 63.67675781
   "001111111010111011", -- Line 1   Column 1528   Coefficient 63.68261719
   "001111111011000001", -- Line 1   Column 1529   Coefficient 63.68847656
   "001111111011000110", -- Line 1   Column 1530   Coefficient 63.69335938
   "001111111011001100", -- Line 1   Column 1531   Coefficient 63.69921875
   "001111111011010010", -- Line 1   Column 1532   Coefficient 63.70507813
   "001111111011011000", -- Line 1   Column 1533   Coefficient 63.71093750
   "001111111011011110", -- Line 1   Column 1534   Coefficient 63.71679688
   "001111111011100011", -- Line 1   Column 1535   Coefficient 63.72167969
   "001111111011101001", -- Line 1   Column 1536   Coefficient 63.72753906
   "001111111011101111", -- Line 1   Column 1537   Coefficient 63.73339844
   "001111111011110101", -- Line 1   Column 1538   Coefficient 63.73925781
   "001111111011111011", -- Line 1   Column 1539   Coefficient 63.74511719
   "001111111100000000", -- Line 1   Column 1540   Coefficient 63.75000000
   "001111111100000110", -- Line 1   Column 1541   Coefficient 63.75585938
   "001111111100001100", -- Line 1   Column 1542   Coefficient 63.76171875
   "001111111100010010", -- Line 1   Column 1543   Coefficient 63.76757813
   "001111111100010111", -- Line 1   Column 1544   Coefficient 63.77246094
   "001111111100011101", -- Line 1   Column 1545   Coefficient 63.77832031
   "001111111100100011", -- Line 1   Column 1546   Coefficient 63.78417969
   "001111111100101001", -- Line 1   Column 1547   Coefficient 63.79003906
   "001111111100101111", -- Line 1   Column 1548   Coefficient 63.79589844
   "001111111100110100", -- Line 1   Column 1549   Coefficient 63.80078125
   "001111111100111010", -- Line 1   Column 1550   Coefficient 63.80664063
   "001111111101000000", -- Line 1   Column 1551   Coefficient 63.81250000
   "001111111101000101", -- Line 1   Column 1552   Coefficient 63.81738281
   "001111111101001011", -- Line 1   Column 1553   Coefficient 63.82324219
   "001111111101010001", -- Line 1   Column 1554   Coefficient 63.82910156
   "001111111101010111", -- Line 1   Column 1555   Coefficient 63.83496094
   "001111111101011100", -- Line 1   Column 1556   Coefficient 63.83984375
   "001111111101100010", -- Line 1   Column 1557   Coefficient 63.84570313
   "001111111101101000", -- Line 1   Column 1558   Coefficient 63.85156250
   "001111111101101101", -- Line 1   Column 1559   Coefficient 63.85644531
   "001111111101110011", -- Line 1   Column 1560   Coefficient 63.86230469
   "001111111101111001", -- Line 1   Column 1561   Coefficient 63.86816406
   "001111111101111111", -- Line 1   Column 1562   Coefficient 63.87402344
   "001111111110000100", -- Line 1   Column 1563   Coefficient 63.87890625
   "001111111110001010", -- Line 1   Column 1564   Coefficient 63.88476563
   "001111111110010000", -- Line 1   Column 1565   Coefficient 63.89062500
   "001111111110010101", -- Line 1   Column 1566   Coefficient 63.89550781
   "001111111110011011", -- Line 1   Column 1567   Coefficient 63.90136719
   "001111111110100001", -- Line 1   Column 1568   Coefficient 63.90722656
   "001111111110100110", -- Line 1   Column 1569   Coefficient 63.91210938
   "001111111110101100", -- Line 1   Column 1570   Coefficient 63.91796875
   "001111111110110010", -- Line 1   Column 1571   Coefficient 63.92382813
   "001111111110110111", -- Line 1   Column 1572   Coefficient 63.92871094
   "001111111110111101", -- Line 1   Column 1573   Coefficient 63.93457031
   "001111111111000011", -- Line 1   Column 1574   Coefficient 63.94042969
   "001111111111001000", -- Line 1   Column 1575   Coefficient 63.94531250
   "001111111111001110", -- Line 1   Column 1576   Coefficient 63.95117188
   "001111111111010100", -- Line 1   Column 1577   Coefficient 63.95703125
   "001111111111011001", -- Line 1   Column 1578   Coefficient 63.96191406
   "001111111111011111", -- Line 1   Column 1579   Coefficient 63.96777344
   "001111111111100100", -- Line 1   Column 1580   Coefficient 63.97265625
   "001111111111101010", -- Line 1   Column 1581   Coefficient 63.97851563
   "001111111111110000", -- Line 1   Column 1582   Coefficient 63.98437500
   "001111111111110101", -- Line 1   Column 1583   Coefficient 63.98925781
   "001111111111111011", -- Line 1   Column 1584   Coefficient 63.99511719
   "010000000000000001", -- Line 1   Column 1585   Coefficient 64.00097656
   "010000000000000110", -- Line 1   Column 1586   Coefficient 64.00585938
   "010000000000001100", -- Line 1   Column 1587   Coefficient 64.01171875
   "010000000000010001", -- Line 1   Column 1588   Coefficient 64.01660156
   "010000000000010111", -- Line 1   Column 1589   Coefficient 64.02246094
   "010000000000011101", -- Line 1   Column 1590   Coefficient 64.02832031
   "010000000000100010", -- Line 1   Column 1591   Coefficient 64.03320313
   "010000000000101000", -- Line 1   Column 1592   Coefficient 64.03906250
   "010000000000101101", -- Line 1   Column 1593   Coefficient 64.04394531
   "010000000000110011", -- Line 1   Column 1594   Coefficient 64.04980469
   "010000000000111001", -- Line 1   Column 1595   Coefficient 64.05566406
   "010000000000111110", -- Line 1   Column 1596   Coefficient 64.06054688
   "010000000001000100", -- Line 1   Column 1597   Coefficient 64.06640625
   "010000000001001001", -- Line 1   Column 1598   Coefficient 64.07128906
   "010000000001001111", -- Line 1   Column 1599   Coefficient 64.07714844
   "010000000001010100", -- Line 1   Column 1600   Coefficient 64.08203125
   "010000000001011010", -- Line 1   Column 1601   Coefficient 64.08789063
   "010000000001011111", -- Line 1   Column 1602   Coefficient 64.09277344
   "010000000001100101", -- Line 1   Column 1603   Coefficient 64.09863281
   "010000000001101011", -- Line 1   Column 1604   Coefficient 64.10449219
   "010000000001110000", -- Line 1   Column 1605   Coefficient 64.10937500
   "010000000001110110", -- Line 1   Column 1606   Coefficient 64.11523438
   "010000000001111011", -- Line 1   Column 1607   Coefficient 64.12011719
   "010000000010000001", -- Line 1   Column 1608   Coefficient 64.12597656
   "010000000010000110", -- Line 1   Column 1609   Coefficient 64.13085938
   "010000000010001100", -- Line 1   Column 1610   Coefficient 64.13671875
   "010000000010010001", -- Line 1   Column 1611   Coefficient 64.14160156
   "010000000010010111", -- Line 1   Column 1612   Coefficient 64.14746094
   "010000000010011100", -- Line 1   Column 1613   Coefficient 64.15234375
   "010000000010100010", -- Line 1   Column 1614   Coefficient 64.15820313
   "010000000010100111", -- Line 1   Column 1615   Coefficient 64.16308594
   "010000000010101101", -- Line 1   Column 1616   Coefficient 64.16894531
   "010000000010110010", -- Line 1   Column 1617   Coefficient 64.17382813
   "010000000010111000", -- Line 1   Column 1618   Coefficient 64.17968750
   "010000000010111101", -- Line 1   Column 1619   Coefficient 64.18457031
   "010000000011000011", -- Line 1   Column 1620   Coefficient 64.19042969
   "010000000011001000", -- Line 1   Column 1621   Coefficient 64.19531250
   "010000000011001110", -- Line 1   Column 1622   Coefficient 64.20117188
   "010000000011010011", -- Line 1   Column 1623   Coefficient 64.20605469
   "010000000011011001", -- Line 1   Column 1624   Coefficient 64.21191406
   "010000000011011110", -- Line 1   Column 1625   Coefficient 64.21679688
   "010000000011100100", -- Line 1   Column 1626   Coefficient 64.22265625
   "010000000011101001", -- Line 1   Column 1627   Coefficient 64.22753906
   "010000000011101111", -- Line 1   Column 1628   Coefficient 64.23339844
   "010000000011110100", -- Line 1   Column 1629   Coefficient 64.23828125
   "010000000011111010", -- Line 1   Column 1630   Coefficient 64.24414063
   "010000000011111111", -- Line 1   Column 1631   Coefficient 64.24902344
   "010000000100000101", -- Line 1   Column 1632   Coefficient 64.25488281
   "010000000100001010", -- Line 1   Column 1633   Coefficient 64.25976563
   "010000000100001111", -- Line 1   Column 1634   Coefficient 64.26464844
   "010000000100010101", -- Line 1   Column 1635   Coefficient 64.27050781
   "010000000100011010", -- Line 1   Column 1636   Coefficient 64.27539063
   "010000000100100000", -- Line 1   Column 1637   Coefficient 64.28125000
   "010000000100100101", -- Line 1   Column 1638   Coefficient 64.28613281
   "010000000100101011", -- Line 1   Column 1639   Coefficient 64.29199219
   "010000000100110000", -- Line 1   Column 1640   Coefficient 64.29687500
   "010000000100110101", -- Line 1   Column 1641   Coefficient 64.30175781
   "010000000100111011", -- Line 1   Column 1642   Coefficient 64.30761719
   "010000000101000000", -- Line 1   Column 1643   Coefficient 64.31250000
   "010000000101000110", -- Line 1   Column 1644   Coefficient 64.31835938
   "010000000101001011", -- Line 1   Column 1645   Coefficient 64.32324219
   "010000000101010000", -- Line 1   Column 1646   Coefficient 64.32812500
   "010000000101010110", -- Line 1   Column 1647   Coefficient 64.33398438
   "010000000101011011", -- Line 1   Column 1648   Coefficient 64.33886719
   "010000000101100001", -- Line 1   Column 1649   Coefficient 64.34472656
   "010000000101100110", -- Line 1   Column 1650   Coefficient 64.34960938
   "010000000101101011", -- Line 1   Column 1651   Coefficient 64.35449219
   "010000000101110001", -- Line 1   Column 1652   Coefficient 64.36035156
   "010000000101110110", -- Line 1   Column 1653   Coefficient 64.36523438
   "010000000101111100", -- Line 1   Column 1654   Coefficient 64.37109375
   "010000000110000001", -- Line 1   Column 1655   Coefficient 64.37597656
   "010000000110000110", -- Line 1   Column 1656   Coefficient 64.38085938
   "010000000110001100", -- Line 1   Column 1657   Coefficient 64.38671875
   "010000000110010001", -- Line 1   Column 1658   Coefficient 64.39160156
   "010000000110010110", -- Line 1   Column 1659   Coefficient 64.39648438
   "010000000110011100", -- Line 1   Column 1660   Coefficient 64.40234375
   "010000000110100001", -- Line 1   Column 1661   Coefficient 64.40722656
   "010000000110100111", -- Line 1   Column 1662   Coefficient 64.41308594
   "010000000110101100", -- Line 1   Column 1663   Coefficient 64.41796875
   "010000000110110001", -- Line 1   Column 1664   Coefficient 64.42285156
   "010000000110110111", -- Line 1   Column 1665   Coefficient 64.42871094
   "010000000110111100", -- Line 1   Column 1666   Coefficient 64.43359375
   "010000000111000001", -- Line 1   Column 1667   Coefficient 64.43847656
   "010000000111000111", -- Line 1   Column 1668   Coefficient 64.44433594
   "010000000111001100", -- Line 1   Column 1669   Coefficient 64.44921875
   "010000000111010001", -- Line 1   Column 1670   Coefficient 64.45410156
   "010000000111010111", -- Line 1   Column 1671   Coefficient 64.45996094
   "010000000111011100", -- Line 1   Column 1672   Coefficient 64.46484375
   "010000000111100001", -- Line 1   Column 1673   Coefficient 64.46972656
   "010000000111100111", -- Line 1   Column 1674   Coefficient 64.47558594
   "010000000111101100", -- Line 1   Column 1675   Coefficient 64.48046875
   "010000000111110001", -- Line 1   Column 1676   Coefficient 64.48535156
   "010000000111110110", -- Line 1   Column 1677   Coefficient 64.49023438
   "010000000111111100", -- Line 1   Column 1678   Coefficient 64.49609375
   "010000001000000001", -- Line 1   Column 1679   Coefficient 64.50097656
   "010000001000000110", -- Line 1   Column 1680   Coefficient 64.50585938
   "010000001000001100", -- Line 1   Column 1681   Coefficient 64.51171875
   "010000001000010001", -- Line 1   Column 1682   Coefficient 64.51660156
   "010000001000010110", -- Line 1   Column 1683   Coefficient 64.52148438
   "010000001000011011", -- Line 1   Column 1684   Coefficient 64.52636719
   "010000001000100001", -- Line 1   Column 1685   Coefficient 64.53222656
   "010000001000100110", -- Line 1   Column 1686   Coefficient 64.53710938
   "010000001000101011", -- Line 1   Column 1687   Coefficient 64.54199219
   "010000001000110001", -- Line 1   Column 1688   Coefficient 64.54785156
   "010000001000110110", -- Line 1   Column 1689   Coefficient 64.55273438
   "010000001000111011", -- Line 1   Column 1690   Coefficient 64.55761719
   "010000001001000000", -- Line 1   Column 1691   Coefficient 64.56250000
   "010000001001000110", -- Line 1   Column 1692   Coefficient 64.56835938
   "010000001001001011", -- Line 1   Column 1693   Coefficient 64.57324219
   "010000001001010000", -- Line 1   Column 1694   Coefficient 64.57812500
   "010000001001010101", -- Line 1   Column 1695   Coefficient 64.58300781
   "010000001001011011", -- Line 1   Column 1696   Coefficient 64.58886719
   "010000001001100000", -- Line 1   Column 1697   Coefficient 64.59375000
   "010000001001100101", -- Line 1   Column 1698   Coefficient 64.59863281
   "010000001001101010", -- Line 1   Column 1699   Coefficient 64.60351563
   "010000001001110000", -- Line 1   Column 1700   Coefficient 64.60937500
   "010000001001110101", -- Line 1   Column 1701   Coefficient 64.61425781
   "010000001001111010", -- Line 1   Column 1702   Coefficient 64.61914063
   "010000001001111111", -- Line 1   Column 1703   Coefficient 64.62402344
   "010000001010000100", -- Line 1   Column 1704   Coefficient 64.62890625
   "010000001010001010", -- Line 1   Column 1705   Coefficient 64.63476563
   "010000001010001111", -- Line 1   Column 1706   Coefficient 64.63964844
   "010000001010010100", -- Line 1   Column 1707   Coefficient 64.64453125
   "010000001010011001", -- Line 1   Column 1708   Coefficient 64.64941406
   "010000001010011111", -- Line 1   Column 1709   Coefficient 64.65527344
   "010000001010100100", -- Line 1   Column 1710   Coefficient 64.66015625
   "010000001010101001", -- Line 1   Column 1711   Coefficient 64.66503906
   "010000001010101110", -- Line 1   Column 1712   Coefficient 64.66992188
   "010000001010110011", -- Line 1   Column 1713   Coefficient 64.67480469
   "010000001010111001", -- Line 1   Column 1714   Coefficient 64.68066406
   "010000001010111110", -- Line 1   Column 1715   Coefficient 64.68554688
   "010000001011000011", -- Line 1   Column 1716   Coefficient 64.69042969
   "010000001011001000", -- Line 1   Column 1717   Coefficient 64.69531250
   "010000001011001101", -- Line 1   Column 1718   Coefficient 64.70019531
   "010000001011010010", -- Line 1   Column 1719   Coefficient 64.70507813
   "010000001011011000", -- Line 1   Column 1720   Coefficient 64.71093750
   "010000001011011101", -- Line 1   Column 1721   Coefficient 64.71582031
   "010000001011100010", -- Line 1   Column 1722   Coefficient 64.72070313
   "010000001011100111", -- Line 1   Column 1723   Coefficient 64.72558594
   "010000001011101100", -- Line 1   Column 1724   Coefficient 64.73046875
   "010000001011110001", -- Line 1   Column 1725   Coefficient 64.73535156
   "010000001011110111", -- Line 1   Column 1726   Coefficient 64.74121094
   "010000001011111100", -- Line 1   Column 1727   Coefficient 64.74609375
   "010000001100000001", -- Line 1   Column 1728   Coefficient 64.75097656
   "010000001100000110", -- Line 1   Column 1729   Coefficient 64.75585938
   "010000001100001011", -- Line 1   Column 1730   Coefficient 64.76074219
   "010000001100010000", -- Line 1   Column 1731   Coefficient 64.76562500
   "010000001100010101", -- Line 1   Column 1732   Coefficient 64.77050781
   "010000001100011011", -- Line 1   Column 1733   Coefficient 64.77636719
   "010000001100100000", -- Line 1   Column 1734   Coefficient 64.78125000
   "010000001100100101", -- Line 1   Column 1735   Coefficient 64.78613281
   "010000001100101010", -- Line 1   Column 1736   Coefficient 64.79101563
   "010000001100101111", -- Line 1   Column 1737   Coefficient 64.79589844
   "010000001100110100", -- Line 1   Column 1738   Coefficient 64.80078125
   "010000001100111001", -- Line 1   Column 1739   Coefficient 64.80566406
   "010000001100111110", -- Line 1   Column 1740   Coefficient 64.81054688
   "010000001101000100", -- Line 1   Column 1741   Coefficient 64.81640625
   "010000001101001001", -- Line 1   Column 1742   Coefficient 64.82128906
   "010000001101001110", -- Line 1   Column 1743   Coefficient 64.82617188
   "010000001101010011", -- Line 1   Column 1744   Coefficient 64.83105469
   "010000001101011000", -- Line 1   Column 1745   Coefficient 64.83593750
   "010000001101011101", -- Line 1   Column 1746   Coefficient 64.84082031
   "010000001101100010", -- Line 1   Column 1747   Coefficient 64.84570313
   "010000001101100111", -- Line 1   Column 1748   Coefficient 64.85058594
   "010000001101101100", -- Line 1   Column 1749   Coefficient 64.85546875
   "010000001101110001", -- Line 1   Column 1750   Coefficient 64.86035156
   "010000001101110111", -- Line 1   Column 1751   Coefficient 64.86621094
   "010000001101111100", -- Line 1   Column 1752   Coefficient 64.87109375
   "010000001110000001", -- Line 1   Column 1753   Coefficient 64.87597656
   "010000001110000110", -- Line 1   Column 1754   Coefficient 64.88085938
   "010000001110001011", -- Line 1   Column 1755   Coefficient 64.88574219
   "010000001110010000", -- Line 1   Column 1756   Coefficient 64.89062500
   "010000001110010101", -- Line 1   Column 1757   Coefficient 64.89550781
   "010000001110011010", -- Line 1   Column 1758   Coefficient 64.90039063
   "010000001110011111", -- Line 1   Column 1759   Coefficient 64.90527344
   "010000001110100100", -- Line 1   Column 1760   Coefficient 64.91015625
   "010000001110101001", -- Line 1   Column 1761   Coefficient 64.91503906
   "010000001110101110", -- Line 1   Column 1762   Coefficient 64.91992188
   "010000001110110011", -- Line 1   Column 1763   Coefficient 64.92480469
   "010000001110111000", -- Line 1   Column 1764   Coefficient 64.92968750
   "010000001110111101", -- Line 1   Column 1765   Coefficient 64.93457031
   "010000001111000010", -- Line 1   Column 1766   Coefficient 64.93945313
   "010000001111000111", -- Line 1   Column 1767   Coefficient 64.94433594
   "010000001111001100", -- Line 1   Column 1768   Coefficient 64.94921875
   "010000001111010001", -- Line 1   Column 1769   Coefficient 64.95410156
   "010000001111010110", -- Line 1   Column 1770   Coefficient 64.95898438
   "010000001111011100", -- Line 1   Column 1771   Coefficient 64.96484375
   "010000001111100001", -- Line 1   Column 1772   Coefficient 64.96972656
   "010000001111100110", -- Line 1   Column 1773   Coefficient 64.97460938
   "010000001111101011", -- Line 1   Column 1774   Coefficient 64.97949219
   "010000001111110000", -- Line 1   Column 1775   Coefficient 64.98437500
   "010000001111110101", -- Line 1   Column 1776   Coefficient 64.98925781
   "010000001111111010", -- Line 1   Column 1777   Coefficient 64.99414063
   "010000001111111111", -- Line 1   Column 1778   Coefficient 64.99902344
   "010000010000000100", -- Line 1   Column 1779   Coefficient 65.00390625
   "010000010000001001", -- Line 1   Column 1780   Coefficient 65.00878906
   "010000010000001110", -- Line 1   Column 1781   Coefficient 65.01367188
   "010000010000010011", -- Line 1   Column 1782   Coefficient 65.01855469
   "010000010000011000", -- Line 1   Column 1783   Coefficient 65.02343750
   "010000010000011101", -- Line 1   Column 1784   Coefficient 65.02832031
   "010000010000100010", -- Line 1   Column 1785   Coefficient 65.03320313
   "010000010000100111", -- Line 1   Column 1786   Coefficient 65.03808594
   "010000010000101100", -- Line 1   Column 1787   Coefficient 65.04296875
   "010000010000110000", -- Line 1   Column 1788   Coefficient 65.04687500
   "010000010000110101", -- Line 1   Column 1789   Coefficient 65.05175781
   "010000010000111010", -- Line 1   Column 1790   Coefficient 65.05664063
   "010000010000111111", -- Line 1   Column 1791   Coefficient 65.06152344
   "010000010001000100", -- Line 1   Column 1792   Coefficient 65.06640625
   "010000010001001001", -- Line 1   Column 1793   Coefficient 65.07128906
   "010000010001001110", -- Line 1   Column 1794   Coefficient 65.07617188
   "010000010001010011", -- Line 1   Column 1795   Coefficient 65.08105469
   "010000010001011000", -- Line 1   Column 1796   Coefficient 65.08593750
   "010000010001011101", -- Line 1   Column 1797   Coefficient 65.09082031
   "010000010001100010", -- Line 1   Column 1798   Coefficient 65.09570313
   "010000010001100111", -- Line 1   Column 1799   Coefficient 65.10058594
   "010000010001101100", -- Line 1   Column 1800   Coefficient 65.10546875
   "010000010001110001", -- Line 1   Column 1801   Coefficient 65.11035156
   "010000010001110110", -- Line 1   Column 1802   Coefficient 65.11523438
   "010000010001111011", -- Line 1   Column 1803   Coefficient 65.12011719
   "010000010010000000", -- Line 1   Column 1804   Coefficient 65.12500000
   "010000010010000101", -- Line 1   Column 1805   Coefficient 65.12988281
   "010000010010001010", -- Line 1   Column 1806   Coefficient 65.13476563
   "010000010010001111", -- Line 1   Column 1807   Coefficient 65.13964844
   "010000010010010011", -- Line 1   Column 1808   Coefficient 65.14355469
   "010000010010011000", -- Line 1   Column 1809   Coefficient 65.14843750
   "010000010010011101", -- Line 1   Column 1810   Coefficient 65.15332031
   "010000010010100010", -- Line 1   Column 1811   Coefficient 65.15820313
   "010000010010100111", -- Line 1   Column 1812   Coefficient 65.16308594
   "010000010010101100", -- Line 1   Column 1813   Coefficient 65.16796875
   "010000010010110001", -- Line 1   Column 1814   Coefficient 65.17285156
   "010000010010110110", -- Line 1   Column 1815   Coefficient 65.17773438
   "010000010010111011", -- Line 1   Column 1816   Coefficient 65.18261719
   "010000010011000000", -- Line 1   Column 1817   Coefficient 65.18750000
   "010000010011000100", -- Line 1   Column 1818   Coefficient 65.19140625
   "010000010011001001", -- Line 1   Column 1819   Coefficient 65.19628906
   "010000010011001110", -- Line 1   Column 1820   Coefficient 65.20117188
   "010000010011010011", -- Line 1   Column 1821   Coefficient 65.20605469
   "010000010011011000", -- Line 1   Column 1822   Coefficient 65.21093750
   "010000010011011101", -- Line 1   Column 1823   Coefficient 65.21582031
   "010000010011100010", -- Line 1   Column 1824   Coefficient 65.22070313
   "010000010011100111", -- Line 1   Column 1825   Coefficient 65.22558594
   "010000010011101100", -- Line 1   Column 1826   Coefficient 65.23046875
   "010000010011110000", -- Line 1   Column 1827   Coefficient 65.23437500
   "010000010011110101", -- Line 1   Column 1828   Coefficient 65.23925781
   "010000010011111010", -- Line 1   Column 1829   Coefficient 65.24414063
   "010000010011111111", -- Line 1   Column 1830   Coefficient 65.24902344
   "010000010100000100", -- Line 1   Column 1831   Coefficient 65.25390625
   "010000010100001001", -- Line 1   Column 1832   Coefficient 65.25878906
   "010000010100001110", -- Line 1   Column 1833   Coefficient 65.26367188
   "010000010100010010", -- Line 1   Column 1834   Coefficient 65.26757813
   "010000010100010111", -- Line 1   Column 1835   Coefficient 65.27246094
   "010000010100011100", -- Line 1   Column 1836   Coefficient 65.27734375
   "010000010100100001", -- Line 1   Column 1837   Coefficient 65.28222656
   "010000010100100110", -- Line 1   Column 1838   Coefficient 65.28710938
   "010000010100101011", -- Line 1   Column 1839   Coefficient 65.29199219
   "010000010100101111", -- Line 1   Column 1840   Coefficient 65.29589844
   "010000010100110100", -- Line 1   Column 1841   Coefficient 65.30078125
   "010000010100111001", -- Line 1   Column 1842   Coefficient 65.30566406
   "010000010100111110", -- Line 1   Column 1843   Coefficient 65.31054688
   "010000010101000011", -- Line 1   Column 1844   Coefficient 65.31542969
   "010000010101001000", -- Line 1   Column 1845   Coefficient 65.32031250
   "010000010101001100", -- Line 1   Column 1846   Coefficient 65.32421875
   "010000010101010001", -- Line 1   Column 1847   Coefficient 65.32910156
   "010000010101010110", -- Line 1   Column 1848   Coefficient 65.33398438
   "010000010101011011", -- Line 1   Column 1849   Coefficient 65.33886719
   "010000010101100000", -- Line 1   Column 1850   Coefficient 65.34375000
   "010000010101100100", -- Line 1   Column 1851   Coefficient 65.34765625
   "010000010101101001", -- Line 1   Column 1852   Coefficient 65.35253906
   "010000010101101110", -- Line 1   Column 1853   Coefficient 65.35742188
   "010000010101110011", -- Line 1   Column 1854   Coefficient 65.36230469
   "010000010101111000", -- Line 1   Column 1855   Coefficient 65.36718750
   "010000010101111100", -- Line 1   Column 1856   Coefficient 65.37109375
   "010000010110000001", -- Line 1   Column 1857   Coefficient 65.37597656
   "010000010110000110", -- Line 1   Column 1858   Coefficient 65.38085938
   "010000010110001011", -- Line 1   Column 1859   Coefficient 65.38574219
   "010000010110010000", -- Line 1   Column 1860   Coefficient 65.39062500
   "010000010110010100", -- Line 1   Column 1861   Coefficient 65.39453125
   "010000010110011001", -- Line 1   Column 1862   Coefficient 65.39941406
   "010000010110011110", -- Line 1   Column 1863   Coefficient 65.40429688
   "010000010110100011", -- Line 1   Column 1864   Coefficient 65.40917969
   "010000010110101000", -- Line 1   Column 1865   Coefficient 65.41406250
   "010000010110101100", -- Line 1   Column 1866   Coefficient 65.41796875
   "010000010110110001", -- Line 1   Column 1867   Coefficient 65.42285156
   "010000010110110110", -- Line 1   Column 1868   Coefficient 65.42773438
   "010000010110111011", -- Line 1   Column 1869   Coefficient 65.43261719
   "010000010110111111", -- Line 1   Column 1870   Coefficient 65.43652344
   "010000010111000100", -- Line 1   Column 1871   Coefficient 65.44140625
   "010000010111001001", -- Line 1   Column 1872   Coefficient 65.44628906
   "010000010111001110", -- Line 1   Column 1873   Coefficient 65.45117188
   "010000010111010010", -- Line 1   Column 1874   Coefficient 65.45507813
   "010000010111010111", -- Line 1   Column 1875   Coefficient 65.45996094
   "010000010111011100", -- Line 1   Column 1876   Coefficient 65.46484375
   "010000010111100001", -- Line 1   Column 1877   Coefficient 65.46972656
   "010000010111100101", -- Line 1   Column 1878   Coefficient 65.47363281
   "010000010111101010", -- Line 1   Column 1879   Coefficient 65.47851563
   "010000010111101111", -- Line 1   Column 1880   Coefficient 65.48339844
   "010000010111110011", -- Line 1   Column 1881   Coefficient 65.48730469
   "010000010111111000", -- Line 1   Column 1882   Coefficient 65.49218750
   "010000010111111101", -- Line 1   Column 1883   Coefficient 65.49707031
   "010000011000000010", -- Line 1   Column 1884   Coefficient 65.50195313
   "010000011000000110", -- Line 1   Column 1885   Coefficient 65.50585938
   "010000011000001011", -- Line 1   Column 1886   Coefficient 65.51074219
   "010000011000010000", -- Line 1   Column 1887   Coefficient 65.51562500
   "010000011000010101", -- Line 1   Column 1888   Coefficient 65.52050781
   "010000011000011001", -- Line 1   Column 1889   Coefficient 65.52441406
   "010000011000011110", -- Line 1   Column 1890   Coefficient 65.52929688
   "010000011000100011", -- Line 1   Column 1891   Coefficient 65.53417969
   "010000011000100111", -- Line 1   Column 1892   Coefficient 65.53808594
   "010000011000101100", -- Line 1   Column 1893   Coefficient 65.54296875
   "010000011000110001", -- Line 1   Column 1894   Coefficient 65.54785156
   "010000011000110101", -- Line 1   Column 1895   Coefficient 65.55175781
   "010000011000111010", -- Line 1   Column 1896   Coefficient 65.55664063
   "010000011000111111", -- Line 1   Column 1897   Coefficient 65.56152344
   "010000011001000100", -- Line 1   Column 1898   Coefficient 65.56640625
   "010000011001001000", -- Line 1   Column 1899   Coefficient 65.57031250
   "010000011001001101", -- Line 1   Column 1900   Coefficient 65.57519531
   "010000011001010010", -- Line 1   Column 1901   Coefficient 65.58007813
   "010000011001010110", -- Line 1   Column 1902   Coefficient 65.58398438
   "010000011001011011", -- Line 1   Column 1903   Coefficient 65.58886719
   "010000011001100000", -- Line 1   Column 1904   Coefficient 65.59375000
   "010000011001100100", -- Line 1   Column 1905   Coefficient 65.59765625
   "010000011001101001", -- Line 1   Column 1906   Coefficient 65.60253906
   "010000011001101110", -- Line 1   Column 1907   Coefficient 65.60742188
   "010000011001110010", -- Line 1   Column 1908   Coefficient 65.61132813
   "010000011001110111", -- Line 1   Column 1909   Coefficient 65.61621094
   "010000011001111100", -- Line 1   Column 1910   Coefficient 65.62109375
   "010000011010000000", -- Line 1   Column 1911   Coefficient 65.62500000
   "010000011010000101", -- Line 1   Column 1912   Coefficient 65.62988281
   "010000011010001010", -- Line 1   Column 1913   Coefficient 65.63476563
   "010000011010001110", -- Line 1   Column 1914   Coefficient 65.63867188
   "010000011010010011", -- Line 1   Column 1915   Coefficient 65.64355469
   "010000011010010111", -- Line 1   Column 1916   Coefficient 65.64746094
   "010000011010011100", -- Line 1   Column 1917   Coefficient 65.65234375
   "010000011010100001", -- Line 1   Column 1918   Coefficient 65.65722656
   "010000011010100101", -- Line 1   Column 1919   Coefficient 65.66113281
   "010000011010101010", -- Line 1   Column 1920   Coefficient 65.66601563
   "010000011010101111", -- Line 1   Column 1921   Coefficient 65.67089844
   "010000011010110011", -- Line 1   Column 1922   Coefficient 65.67480469
   "010000011010111000", -- Line 1   Column 1923   Coefficient 65.67968750
   "010000011010111101", -- Line 1   Column 1924   Coefficient 65.68457031
   "010000011011000001", -- Line 1   Column 1925   Coefficient 65.68847656
   "010000011011000110", -- Line 1   Column 1926   Coefficient 65.69335938
   "010000011011001010", -- Line 1   Column 1927   Coefficient 65.69726563
   "010000011011001111", -- Line 1   Column 1928   Coefficient 65.70214844
   "010000011011010100", -- Line 1   Column 1929   Coefficient 65.70703125
   "010000011011011000", -- Line 1   Column 1930   Coefficient 65.71093750
   "010000011011011101", -- Line 1   Column 1931   Coefficient 65.71582031
   "010000011011100001", -- Line 1   Column 1932   Coefficient 65.71972656
   "010000011011100110", -- Line 1   Column 1933   Coefficient 65.72460938
   "010000011011101011", -- Line 1   Column 1934   Coefficient 65.72949219
   "010000011011101111", -- Line 1   Column 1935   Coefficient 65.73339844
   "010000011011110100", -- Line 1   Column 1936   Coefficient 65.73828125
   "010000011011111000", -- Line 1   Column 1937   Coefficient 65.74218750
   "010000011011111101", -- Line 1   Column 1938   Coefficient 65.74707031
   "010000011100000010", -- Line 1   Column 1939   Coefficient 65.75195313
   "010000011100000110", -- Line 1   Column 1940   Coefficient 65.75585938
   "010000011100001011", -- Line 1   Column 1941   Coefficient 65.76074219
   "010000011100001111", -- Line 1   Column 1942   Coefficient 65.76464844
   "010000011100010100", -- Line 1   Column 1943   Coefficient 65.76953125
   "010000011100011000", -- Line 1   Column 1944   Coefficient 65.77343750
   "010000011100011101", -- Line 1   Column 1945   Coefficient 65.77832031
   "010000011100100010", -- Line 1   Column 1946   Coefficient 65.78320313
   "010000011100100110", -- Line 1   Column 1947   Coefficient 65.78710938
   "010000011100101011", -- Line 1   Column 1948   Coefficient 65.79199219
   "010000011100101111", -- Line 1   Column 1949   Coefficient 65.79589844
   "010000011100110100", -- Line 1   Column 1950   Coefficient 65.80078125
   "010000011100111000", -- Line 1   Column 1951   Coefficient 65.80468750
   "010000011100111101", -- Line 1   Column 1952   Coefficient 65.80957031
   "010000011101000010", -- Line 1   Column 1953   Coefficient 65.81445313
   "010000011101000110", -- Line 1   Column 1954   Coefficient 65.81835938
   "010000011101001011", -- Line 1   Column 1955   Coefficient 65.82324219
   "010000011101001111", -- Line 1   Column 1956   Coefficient 65.82714844
   "010000011101010100", -- Line 1   Column 1957   Coefficient 65.83203125
   "010000011101011000", -- Line 1   Column 1958   Coefficient 65.83593750
   "010000011101011101", -- Line 1   Column 1959   Coefficient 65.84082031
   "010000011101100001", -- Line 1   Column 1960   Coefficient 65.84472656
   "010000011101100110", -- Line 1   Column 1961   Coefficient 65.84960938
   "010000011101101010", -- Line 1   Column 1962   Coefficient 65.85351563
   "010000011101101111", -- Line 1   Column 1963   Coefficient 65.85839844
   "010000011101110100", -- Line 1   Column 1964   Coefficient 65.86328125
   "010000011101111000", -- Line 1   Column 1965   Coefficient 65.86718750
   "010000011101111101", -- Line 1   Column 1966   Coefficient 65.87207031
   "010000011110000001", -- Line 1   Column 1967   Coefficient 65.87597656
   "010000011110000110", -- Line 1   Column 1968   Coefficient 65.88085938
   "010000011110001010", -- Line 1   Column 1969   Coefficient 65.88476563
   "010000011110001111", -- Line 1   Column 1970   Coefficient 65.88964844
   "010000011110010011", -- Line 1   Column 1971   Coefficient 65.89355469
   "010000011110011000", -- Line 1   Column 1972   Coefficient 65.89843750
   "010000011110011100", -- Line 1   Column 1973   Coefficient 65.90234375
   "010000011110100001", -- Line 1   Column 1974   Coefficient 65.90722656
   "010000011110100101", -- Line 1   Column 1975   Coefficient 65.91113281
   "010000011110101010", -- Line 1   Column 1976   Coefficient 65.91601563
   "010000011110101110", -- Line 1   Column 1977   Coefficient 65.91992188
   "010000011110110011", -- Line 1   Column 1978   Coefficient 65.92480469
   "010000011110110111", -- Line 1   Column 1979   Coefficient 65.92871094
   "010000011110111100", -- Line 1   Column 1980   Coefficient 65.93359375
   "010000011111000000", -- Line 1   Column 1981   Coefficient 65.93750000
   "010000011111000101", -- Line 1   Column 1982   Coefficient 65.94238281
   "010000011111001001", -- Line 1   Column 1983   Coefficient 65.94628906
   "010000011111001110", -- Line 1   Column 1984   Coefficient 65.95117188
   "010000011111010010", -- Line 1   Column 1985   Coefficient 65.95507813
   "010000011111010111", -- Line 1   Column 1986   Coefficient 65.95996094
   "010000011111011011", -- Line 1   Column 1987   Coefficient 65.96386719
   "010000011111100000", -- Line 1   Column 1988   Coefficient 65.96875000
   "010000011111100100", -- Line 1   Column 1989   Coefficient 65.97265625
   "010000011111101001", -- Line 1   Column 1990   Coefficient 65.97753906
   "010000011111101101", -- Line 1   Column 1991   Coefficient 65.98144531
   "010000011111110001", -- Line 1   Column 1992   Coefficient 65.98535156
   "010000011111110110", -- Line 1   Column 1993   Coefficient 65.99023438
   "010000011111111010", -- Line 1   Column 1994   Coefficient 65.99414063
   "010000011111111111", -- Line 1   Column 1995   Coefficient 65.99902344
   "010000100000000011", -- Line 1   Column 1996   Coefficient 66.00292969
   "010000100000001000", -- Line 1   Column 1997   Coefficient 66.00781250
   "010000100000001100", -- Line 1   Column 1998   Coefficient 66.01171875
   "010000100000010001", -- Line 1   Column 1999   Coefficient 66.01660156
   "010000100000010101", -- Line 1   Column 2000   Coefficient 66.02050781
   "010000100000011010", -- Line 1   Column 2001   Coefficient 66.02539063
   "010000100000011110", -- Line 1   Column 2002   Coefficient 66.02929688
   "010000100000100010", -- Line 1   Column 2003   Coefficient 66.03320313
   "010000100000100111", -- Line 1   Column 2004   Coefficient 66.03808594
   "010000100000101011", -- Line 1   Column 2005   Coefficient 66.04199219
   "010000100000110000", -- Line 1   Column 2006   Coefficient 66.04687500
   "010000100000110100", -- Line 1   Column 2007   Coefficient 66.05078125
   "010000100000111001", -- Line 1   Column 2008   Coefficient 66.05566406
   "010000100000111101", -- Line 1   Column 2009   Coefficient 66.05957031
   "010000100001000001", -- Line 1   Column 2010   Coefficient 66.06347656
   "010000100001000110", -- Line 1   Column 2011   Coefficient 66.06835938
   "010000100001001010", -- Line 1   Column 2012   Coefficient 66.07226563
   "010000100001001111", -- Line 1   Column 2013   Coefficient 66.07714844
   "010000100001010011", -- Line 1   Column 2014   Coefficient 66.08105469
   "010000100001011000", -- Line 1   Column 2015   Coefficient 66.08593750
   "010000100001011100", -- Line 1   Column 2016   Coefficient 66.08984375
   "010000100001100000", -- Line 1   Column 2017   Coefficient 66.09375000
   "010000100001100101", -- Line 1   Column 2018   Coefficient 66.09863281
   "010000100001101001", -- Line 1   Column 2019   Coefficient 66.10253906
   "010000100001101110", -- Line 1   Column 2020   Coefficient 66.10742188
   "010000100001110010", -- Line 1   Column 2021   Coefficient 66.11132813
   "010000100001110110", -- Line 1   Column 2022   Coefficient 66.11523438
   "010000100001111011", -- Line 1   Column 2023   Coefficient 66.12011719
   "010000100001111111", -- Line 1   Column 2024   Coefficient 66.12402344
   "010000100010000100", -- Line 1   Column 2025   Coefficient 66.12890625
   "010000100010001000", -- Line 1   Column 2026   Coefficient 66.13281250
   "010000100010001100", -- Line 1   Column 2027   Coefficient 66.13671875
   "010000100010010001", -- Line 1   Column 2028   Coefficient 66.14160156
   "010000100010010101", -- Line 1   Column 2029   Coefficient 66.14550781
   "010000100010011010", -- Line 1   Column 2030   Coefficient 66.15039063
   "010000100010011110", -- Line 1   Column 2031   Coefficient 66.15429688
   "010000100010100010", -- Line 1   Column 2032   Coefficient 66.15820313
   "010000100010100111", -- Line 1   Column 2033   Coefficient 66.16308594
   "010000100010101011", -- Line 1   Column 2034   Coefficient 66.16699219
   "010000100010101111", -- Line 1   Column 2035   Coefficient 66.17089844
   "010000100010110100", -- Line 1   Column 2036   Coefficient 66.17578125
   "010000100010111000", -- Line 1   Column 2037   Coefficient 66.17968750
   "010000100010111101", -- Line 1   Column 2038   Coefficient 66.18457031
   "010000100011000001", -- Line 1   Column 2039   Coefficient 66.18847656
   "010000100011000101", -- Line 1   Column 2040   Coefficient 66.19238281
   "010000100011001010", -- Line 1   Column 2041   Coefficient 66.19726563
   "010000100011001110", -- Line 1   Column 2042   Coefficient 66.20117188
   "010000100011010010", -- Line 1   Column 2043   Coefficient 66.20507813
   "010000100011010111", -- Line 1   Column 2044   Coefficient 66.20996094
   "010000100011011011", -- Line 1   Column 2045   Coefficient 66.21386719
   "010000100011011111", -- Line 1   Column 2046   Coefficient 66.21777344
   "010000100011100100", -- Line 1   Column 2047   Coefficient 66.22265625
   "010000100011101000", -- Line 1   Column 2048   Coefficient 66.22656250
   "010000100011101100", -- Line 1   Column 2049   Coefficient 66.23046875
   "010000100011110001", -- Line 1   Column 2050   Coefficient 66.23535156
   "010000100011110101", -- Line 1   Column 2051   Coefficient 66.23925781
   "010000100011111001", -- Line 1   Column 2052   Coefficient 66.24316406
   "010000100011111110", -- Line 1   Column 2053   Coefficient 66.24804688
   "010000100100000010", -- Line 1   Column 2054   Coefficient 66.25195313
   "010000100100000110", -- Line 1   Column 2055   Coefficient 66.25585938
   "010000100100001011", -- Line 1   Column 2056   Coefficient 66.26074219
   "010000100100001111", -- Line 1   Column 2057   Coefficient 66.26464844
   "010000100100010011", -- Line 1   Column 2058   Coefficient 66.26855469
   "010000100100011000", -- Line 1   Column 2059   Coefficient 66.27343750
   "010000100100011100", -- Line 1   Column 2060   Coefficient 66.27734375
   "010000100100100000", -- Line 1   Column 2061   Coefficient 66.28125000
   "010000100100100101", -- Line 1   Column 2062   Coefficient 66.28613281
   "010000100100101001", -- Line 1   Column 2063   Coefficient 66.29003906
   "010000100100101101", -- Line 1   Column 2064   Coefficient 66.29394531
   "010000100100110010", -- Line 1   Column 2065   Coefficient 66.29882813
   "010000100100110110", -- Line 1   Column 2066   Coefficient 66.30273438
   "010000100100111010", -- Line 1   Column 2067   Coefficient 66.30664063
   "010000100100111110", -- Line 1   Column 2068   Coefficient 66.31054688
   "010000100101000011", -- Line 1   Column 2069   Coefficient 66.31542969
   "010000100101000111", -- Line 1   Column 2070   Coefficient 66.31933594
   "010000100101001011", -- Line 1   Column 2071   Coefficient 66.32324219
   "010000100101010000", -- Line 1   Column 2072   Coefficient 66.32812500
   "010000100101010100", -- Line 1   Column 2073   Coefficient 66.33203125
   "010000100101011000", -- Line 1   Column 2074   Coefficient 66.33593750
   "010000100101011101", -- Line 1   Column 2075   Coefficient 66.34082031
   "010000100101100001", -- Line 1   Column 2076   Coefficient 66.34472656
   "010000100101100101", -- Line 1   Column 2077   Coefficient 66.34863281
   "010000100101101001", -- Line 1   Column 2078   Coefficient 66.35253906
   "010000100101101110", -- Line 1   Column 2079   Coefficient 66.35742188
   "010000100101110010", -- Line 1   Column 2080   Coefficient 66.36132813
   "010000100101110110", -- Line 1   Column 2081   Coefficient 66.36523438
   "010000100101111010", -- Line 1   Column 2082   Coefficient 66.36914063
   "010000100101111111", -- Line 1   Column 2083   Coefficient 66.37402344
   "010000100110000011", -- Line 1   Column 2084   Coefficient 66.37792969
   "010000100110000111", -- Line 1   Column 2085   Coefficient 66.38183594
   "010000100110001100", -- Line 1   Column 2086   Coefficient 66.38671875
   "010000100110010000", -- Line 1   Column 2087   Coefficient 66.39062500
   "010000100110010100", -- Line 1   Column 2088   Coefficient 66.39453125
   "010000100110011000", -- Line 1   Column 2089   Coefficient 66.39843750
   "010000100110011101", -- Line 1   Column 2090   Coefficient 66.40332031
   "010000100110100001", -- Line 1   Column 2091   Coefficient 66.40722656
   "010000100110100101", -- Line 1   Column 2092   Coefficient 66.41113281
   "010000100110101001", -- Line 1   Column 2093   Coefficient 66.41503906
   "010000100110101110", -- Line 1   Column 2094   Coefficient 66.41992188
   "010000100110110010", -- Line 1   Column 2095   Coefficient 66.42382813
   "010000100110110110", -- Line 1   Column 2096   Coefficient 66.42773438
   "010000100110111010", -- Line 1   Column 2097   Coefficient 66.43164063
   "010000100110111111", -- Line 1   Column 2098   Coefficient 66.43652344
   "010000100111000011", -- Line 1   Column 2099   Coefficient 66.44042969
   "010000100111000111", -- Line 1   Column 2100   Coefficient 66.44433594
   "010000100111001011", -- Line 1   Column 2101   Coefficient 66.44824219
   "010000100111010000", -- Line 1   Column 2102   Coefficient 66.45312500
   "010000100111010100", -- Line 1   Column 2103   Coefficient 66.45703125
   "010000100111011000", -- Line 1   Column 2104   Coefficient 66.46093750
   "010000100111011100", -- Line 1   Column 2105   Coefficient 66.46484375
   "010000100111100000", -- Line 1   Column 2106   Coefficient 66.46875000
   "010000100111100101", -- Line 1   Column 2107   Coefficient 66.47363281
   "010000100111101001", -- Line 1   Column 2108   Coefficient 66.47753906
   "010000100111101101", -- Line 1   Column 2109   Coefficient 66.48144531
   "010000100111110001", -- Line 1   Column 2110   Coefficient 66.48535156
   "010000100111110110", -- Line 1   Column 2111   Coefficient 66.49023438
   "010000100111111010", -- Line 1   Column 2112   Coefficient 66.49414063
   "010000100111111110", -- Line 1   Column 2113   Coefficient 66.49804688
   "010000101000000010", -- Line 1   Column 2114   Coefficient 66.50195313
   "010000101000000110", -- Line 1   Column 2115   Coefficient 66.50585938
   "010000101000001011", -- Line 1   Column 2116   Coefficient 66.51074219
   "010000101000001111", -- Line 1   Column 2117   Coefficient 66.51464844
   "010000101000010011", -- Line 1   Column 2118   Coefficient 66.51855469
   "010000101000010111", -- Line 1   Column 2119   Coefficient 66.52246094
   "010000101000011011", -- Line 1   Column 2120   Coefficient 66.52636719
   "010000101000100000", -- Line 1   Column 2121   Coefficient 66.53125000
   "010000101000100100", -- Line 1   Column 2122   Coefficient 66.53515625
   "010000101000101000", -- Line 1   Column 2123   Coefficient 66.53906250
   "010000101000101100", -- Line 1   Column 2124   Coefficient 66.54296875
   "010000101000110000", -- Line 1   Column 2125   Coefficient 66.54687500
   "010000101000110100", -- Line 1   Column 2126   Coefficient 66.55078125
   "010000101000111001", -- Line 1   Column 2127   Coefficient 66.55566406
   "010000101000111101", -- Line 1   Column 2128   Coefficient 66.55957031
   "010000101001000001", -- Line 1   Column 2129   Coefficient 66.56347656
   "010000101001000101", -- Line 1   Column 2130   Coefficient 66.56738281
   "010000101001001001", -- Line 1   Column 2131   Coefficient 66.57128906
   "010000101001001110", -- Line 1   Column 2132   Coefficient 66.57617188
   "010000101001010010", -- Line 1   Column 2133   Coefficient 66.58007813
   "010000101001010110", -- Line 1   Column 2134   Coefficient 66.58398438
   "010000101001011010", -- Line 1   Column 2135   Coefficient 66.58789063
   "010000101001011110", -- Line 1   Column 2136   Coefficient 66.59179688
   "010000101001100010", -- Line 1   Column 2137   Coefficient 66.59570313
   "010000101001100111", -- Line 1   Column 2138   Coefficient 66.60058594
   "010000101001101011", -- Line 1   Column 2139   Coefficient 66.60449219
   "010000101001101111", -- Line 1   Column 2140   Coefficient 66.60839844
   "010000101001110011", -- Line 1   Column 2141   Coefficient 66.61230469
   "010000101001110111", -- Line 1   Column 2142   Coefficient 66.61621094
   "010000101001111011", -- Line 1   Column 2143   Coefficient 66.62011719
   "010000101001111111", -- Line 1   Column 2144   Coefficient 66.62402344
   "010000101010000100", -- Line 1   Column 2145   Coefficient 66.62890625
   "010000101010001000", -- Line 1   Column 2146   Coefficient 66.63281250
   "010000101010001100", -- Line 1   Column 2147   Coefficient 66.63671875
   "010000101010010000", -- Line 1   Column 2148   Coefficient 66.64062500
   "010000101010010100", -- Line 1   Column 2149   Coefficient 66.64453125
   "010000101010011000", -- Line 1   Column 2150   Coefficient 66.64843750
   "010000101010011100", -- Line 1   Column 2151   Coefficient 66.65234375
   "010000101010100001", -- Line 1   Column 2152   Coefficient 66.65722656
   "010000101010100101", -- Line 1   Column 2153   Coefficient 66.66113281
   "010000101010101001", -- Line 1   Column 2154   Coefficient 66.66503906
   "010000101010101101", -- Line 1   Column 2155   Coefficient 66.66894531
   "010000101010110001", -- Line 1   Column 2156   Coefficient 66.67285156
   "010000101010110101", -- Line 1   Column 2157   Coefficient 66.67675781
   "010000101010111001", -- Line 1   Column 2158   Coefficient 66.68066406
   "010000101010111101", -- Line 1   Column 2159   Coefficient 66.68457031
   "010000101011000010", -- Line 1   Column 2160   Coefficient 66.68945313
   "010000101011000110", -- Line 1   Column 2161   Coefficient 66.69335938
   "010000101011001010", -- Line 1   Column 2162   Coefficient 66.69726563
   "010000101011001110", -- Line 1   Column 2163   Coefficient 66.70117188
   "010000101011010010", -- Line 1   Column 2164   Coefficient 66.70507813
   "010000101011010110", -- Line 1   Column 2165   Coefficient 66.70898438
   "010000101011011010", -- Line 1   Column 2166   Coefficient 66.71289063
   "010000101011011110", -- Line 1   Column 2167   Coefficient 66.71679688
   "010000101011100010", -- Line 1   Column 2168   Coefficient 66.72070313
   "010000101011100111", -- Line 1   Column 2169   Coefficient 66.72558594
   "010000101011101011", -- Line 1   Column 2170   Coefficient 66.72949219
   "010000101011101111", -- Line 1   Column 2171   Coefficient 66.73339844
   "010000101011110011", -- Line 1   Column 2172   Coefficient 66.73730469
   "010000101011110111", -- Line 1   Column 2173   Coefficient 66.74121094
   "010000101011111011", -- Line 1   Column 2174   Coefficient 66.74511719
   "010000101011111111", -- Line 1   Column 2175   Coefficient 66.74902344
   "010000101100000011", -- Line 1   Column 2176   Coefficient 66.75292969
   "010000101100000111", -- Line 1   Column 2177   Coefficient 66.75683594
   "010000101100001011", -- Line 1   Column 2178   Coefficient 66.76074219
   "010000101100010000", -- Line 1   Column 2179   Coefficient 66.76562500
   "010000101100010100", -- Line 1   Column 2180   Coefficient 66.76953125
   "010000101100011000", -- Line 1   Column 2181   Coefficient 66.77343750
   "010000101100011100", -- Line 1   Column 2182   Coefficient 66.77734375
   "010000101100100000", -- Line 1   Column 2183   Coefficient 66.78125000
   "010000101100100100", -- Line 1   Column 2184   Coefficient 66.78515625
   "010000101100101000", -- Line 1   Column 2185   Coefficient 66.78906250
   "010000101100101100", -- Line 1   Column 2186   Coefficient 66.79296875
   "010000101100110000", -- Line 1   Column 2187   Coefficient 66.79687500
   "010000101100110100", -- Line 1   Column 2188   Coefficient 66.80078125
   "010000101100111000", -- Line 1   Column 2189   Coefficient 66.80468750
   "010000101100111100", -- Line 1   Column 2190   Coefficient 66.80859375
   "010000101101000000", -- Line 1   Column 2191   Coefficient 66.81250000
   "010000101101000100", -- Line 1   Column 2192   Coefficient 66.81640625
   "010000101101001000", -- Line 1   Column 2193   Coefficient 66.82031250
   "010000101101001101", -- Line 1   Column 2194   Coefficient 66.82519531
   "010000101101010001", -- Line 1   Column 2195   Coefficient 66.82910156
   "010000101101010101", -- Line 1   Column 2196   Coefficient 66.83300781
   "010000101101011001", -- Line 1   Column 2197   Coefficient 66.83691406
   "010000101101011101", -- Line 1   Column 2198   Coefficient 66.84082031
   "010000101101100001", -- Line 1   Column 2199   Coefficient 66.84472656
   "010000101101100101", -- Line 1   Column 2200   Coefficient 66.84863281
   "010000101101101001", -- Line 1   Column 2201   Coefficient 66.85253906
   "010000101101101101", -- Line 1   Column 2202   Coefficient 66.85644531
   "010000101101110001", -- Line 1   Column 2203   Coefficient 66.86035156
   "010000101101110101", -- Line 1   Column 2204   Coefficient 66.86425781
   "010000101101111001", -- Line 1   Column 2205   Coefficient 66.86816406
   "010000101101111101", -- Line 1   Column 2206   Coefficient 66.87207031
   "010000101110000001", -- Line 1   Column 2207   Coefficient 66.87597656
   "010000101110000101", -- Line 1   Column 2208   Coefficient 66.87988281
   "010000101110001001", -- Line 1   Column 2209   Coefficient 66.88378906
   "010000101110001101", -- Line 1   Column 2210   Coefficient 66.88769531
   "010000101110010001", -- Line 1   Column 2211   Coefficient 66.89160156
   "010000101110010101", -- Line 1   Column 2212   Coefficient 66.89550781
   "010000101110011001", -- Line 1   Column 2213   Coefficient 66.89941406
   "010000101110011101", -- Line 1   Column 2214   Coefficient 66.90332031
   "010000101110100001", -- Line 1   Column 2215   Coefficient 66.90722656
   "010000101110100101", -- Line 1   Column 2216   Coefficient 66.91113281
   "010000101110101001", -- Line 1   Column 2217   Coefficient 66.91503906
   "010000101110101101", -- Line 1   Column 2218   Coefficient 66.91894531
   "010000101110110001", -- Line 1   Column 2219   Coefficient 66.92285156
   "010000101110110101", -- Line 1   Column 2220   Coefficient 66.92675781
   "010000101110111001", -- Line 1   Column 2221   Coefficient 66.93066406
   "010000101110111101", -- Line 1   Column 2222   Coefficient 66.93457031
   "010000101111000001", -- Line 1   Column 2223   Coefficient 66.93847656
   "010000101111000101", -- Line 1   Column 2224   Coefficient 66.94238281
   "010000101111001001", -- Line 1   Column 2225   Coefficient 66.94628906
   "010000101111001101", -- Line 1   Column 2226   Coefficient 66.95019531
   "010000101111010001", -- Line 1   Column 2227   Coefficient 66.95410156
   "010000101111010101", -- Line 1   Column 2228   Coefficient 66.95800781
   "010000101111011001", -- Line 1   Column 2229   Coefficient 66.96191406
   "010000101111011101", -- Line 1   Column 2230   Coefficient 66.96582031
   "010000101111100001", -- Line 1   Column 2231   Coefficient 66.96972656
   "010000101111100101", -- Line 1   Column 2232   Coefficient 66.97363281
   "010000101111101001", -- Line 1   Column 2233   Coefficient 66.97753906
   "010000101111101101", -- Line 1   Column 2234   Coefficient 66.98144531
   "010000101111110001", -- Line 1   Column 2235   Coefficient 66.98535156
   "010000101111110101", -- Line 1   Column 2236   Coefficient 66.98925781
   "010000101111111001", -- Line 1   Column 2237   Coefficient 66.99316406
   "010000101111111101", -- Line 1   Column 2238   Coefficient 66.99707031
   "010000110000000001", -- Line 1   Column 2239   Coefficient 67.00097656
   "010000110000000101", -- Line 1   Column 2240   Coefficient 67.00488281
   "010000110000001001", -- Line 1   Column 2241   Coefficient 67.00878906
   "010000110000001101", -- Line 1   Column 2242   Coefficient 67.01269531
   "010000110000010001", -- Line 1   Column 2243   Coefficient 67.01660156
   "010000110000010101", -- Line 1   Column 2244   Coefficient 67.02050781
   "010000110000011001", -- Line 1   Column 2245   Coefficient 67.02441406
   "010000110000011101", -- Line 1   Column 2246   Coefficient 67.02832031
   "010000110000100001", -- Line 1   Column 2247   Coefficient 67.03222656
   "010000110000100101", -- Line 1   Column 2248   Coefficient 67.03613281
   "010000110000101001", -- Line 1   Column 2249   Coefficient 67.04003906
   "010000110000101101", -- Line 1   Column 2250   Coefficient 67.04394531
   "010000110000110001", -- Line 1   Column 2251   Coefficient 67.04785156
   "010000110000110101", -- Line 1   Column 2252   Coefficient 67.05175781
   "010000110000111001", -- Line 1   Column 2253   Coefficient 67.05566406
   "010000110000111100", -- Line 1   Column 2254   Coefficient 67.05859375
   "010000110001000000", -- Line 1   Column 2255   Coefficient 67.06250000
   "010000110001000100", -- Line 1   Column 2256   Coefficient 67.06640625
   "010000110001001000", -- Line 1   Column 2257   Coefficient 67.07031250
   "010000110001001100", -- Line 1   Column 2258   Coefficient 67.07421875
   "010000110001010000", -- Line 1   Column 2259   Coefficient 67.07812500
   "010000110001010100", -- Line 1   Column 2260   Coefficient 67.08203125
   "010000110001011000", -- Line 1   Column 2261   Coefficient 67.08593750
   "010000110001011100", -- Line 1   Column 2262   Coefficient 67.08984375
   "010000110001100000", -- Line 1   Column 2263   Coefficient 67.09375000
   "010000110001100100", -- Line 1   Column 2264   Coefficient 67.09765625
   "010000110001101000", -- Line 1   Column 2265   Coefficient 67.10156250
   "010000110001101100", -- Line 1   Column 2266   Coefficient 67.10546875
   "010000110001110000", -- Line 1   Column 2267   Coefficient 67.10937500
   "010000110001110100", -- Line 1   Column 2268   Coefficient 67.11328125
   "010000110001110111", -- Line 1   Column 2269   Coefficient 67.11621094
   "010000110001111011", -- Line 1   Column 2270   Coefficient 67.12011719
   "010000110001111111", -- Line 1   Column 2271   Coefficient 67.12402344
   "010000110010000011", -- Line 1   Column 2272   Coefficient 67.12792969
   "010000110010000111", -- Line 1   Column 2273   Coefficient 67.13183594
   "010000110010001011", -- Line 1   Column 2274   Coefficient 67.13574219
   "010000110010001111", -- Line 1   Column 2275   Coefficient 67.13964844
   "010000110010010011", -- Line 1   Column 2276   Coefficient 67.14355469
   "010000110010010111", -- Line 1   Column 2277   Coefficient 67.14746094
   "010000110010011011", -- Line 1   Column 2278   Coefficient 67.15136719
   "010000110010011111", -- Line 1   Column 2279   Coefficient 67.15527344
   "010000110010100011", -- Line 1   Column 2280   Coefficient 67.15917969
   "010000110010100110", -- Line 1   Column 2281   Coefficient 67.16210938
   "010000110010101010", -- Line 1   Column 2282   Coefficient 67.16601563
   "010000110010101110", -- Line 1   Column 2283   Coefficient 67.16992188
   "010000110010110010", -- Line 1   Column 2284   Coefficient 67.17382813
   "010000110010110110", -- Line 1   Column 2285   Coefficient 67.17773438
   "010000110010111010", -- Line 1   Column 2286   Coefficient 67.18164063
   "010000110010111110", -- Line 1   Column 2287   Coefficient 67.18554688
   "010000110011000010", -- Line 1   Column 2288   Coefficient 67.18945313
   "010000110011000110", -- Line 1   Column 2289   Coefficient 67.19335938
   "010000110011001001", -- Line 1   Column 2290   Coefficient 67.19628906
   "010000110011001101", -- Line 1   Column 2291   Coefficient 67.20019531
   "010000110011010001", -- Line 1   Column 2292   Coefficient 67.20410156
   "010000110011010101", -- Line 1   Column 2293   Coefficient 67.20800781
   "010000110011011001", -- Line 1   Column 2294   Coefficient 67.21191406
   "010000110011011101", -- Line 1   Column 2295   Coefficient 67.21582031
   "010000110011100001", -- Line 1   Column 2296   Coefficient 67.21972656
   "010000110011100101", -- Line 1   Column 2297   Coefficient 67.22363281
   "010000110011101000", -- Line 1   Column 2298   Coefficient 67.22656250
   "010000110011101100", -- Line 1   Column 2299   Coefficient 67.23046875
   "010000110011110000", -- Line 1   Column 2300   Coefficient 67.23437500
   "010000110011110100", -- Line 1   Column 2301   Coefficient 67.23828125
   "010000110011111000", -- Line 1   Column 2302   Coefficient 67.24218750
   "010000110011111100", -- Line 1   Column 2303   Coefficient 67.24609375
   "010000110100000000", -- Line 1   Column 2304   Coefficient 67.25000000
   "010000110100000100", -- Line 1   Column 2305   Coefficient 67.25390625
   "010000110100000111", -- Line 1   Column 2306   Coefficient 67.25683594
   "010000110100001011", -- Line 1   Column 2307   Coefficient 67.26074219
   "010000110100001111", -- Line 1   Column 2308   Coefficient 67.26464844
   "010000110100010011", -- Line 1   Column 2309   Coefficient 67.26855469
   "010000110100010111", -- Line 1   Column 2310   Coefficient 67.27246094
   "010000110100011011", -- Line 1   Column 2311   Coefficient 67.27636719
   "010000110100011110", -- Line 1   Column 2312   Coefficient 67.27929688
   "010000110100100010", -- Line 1   Column 2313   Coefficient 67.28320313
   "010000110100100110", -- Line 1   Column 2314   Coefficient 67.28710938
   "010000110100101010", -- Line 1   Column 2315   Coefficient 67.29101563
   "010000110100101110", -- Line 1   Column 2316   Coefficient 67.29492188
   "010000110100110010", -- Line 1   Column 2317   Coefficient 67.29882813
   "010000110100110110", -- Line 1   Column 2318   Coefficient 67.30273438
   "010000110100111001", -- Line 1   Column 2319   Coefficient 67.30566406
   "010000110100111101", -- Line 1   Column 2320   Coefficient 67.30957031
   "010000110101000001", -- Line 1   Column 2321   Coefficient 67.31347656
   "010000110101000101", -- Line 1   Column 2322   Coefficient 67.31738281
   "010000110101001001", -- Line 1   Column 2323   Coefficient 67.32128906
   "010000110101001101", -- Line 1   Column 2324   Coefficient 67.32519531
   "010000110101010000", -- Line 1   Column 2325   Coefficient 67.32812500
   "010000110101010100", -- Line 1   Column 2326   Coefficient 67.33203125
   "010000110101011000", -- Line 1   Column 2327   Coefficient 67.33593750
   "010000110101011100", -- Line 1   Column 2328   Coefficient 67.33984375
   "010000110101100000", -- Line 1   Column 2329   Coefficient 67.34375000
   "010000110101100011", -- Line 1   Column 2330   Coefficient 67.34667969
   "010000110101100111", -- Line 1   Column 2331   Coefficient 67.35058594
   "010000110101101011", -- Line 1   Column 2332   Coefficient 67.35449219
   "010000110101101111", -- Line 1   Column 2333   Coefficient 67.35839844
   "010000110101110011", -- Line 1   Column 2334   Coefficient 67.36230469
   "010000110101110111", -- Line 1   Column 2335   Coefficient 67.36621094
   "010000110101111010", -- Line 1   Column 2336   Coefficient 67.36914063
   "010000110101111110", -- Line 1   Column 2337   Coefficient 67.37304688
   "010000110110000010", -- Line 1   Column 2338   Coefficient 67.37695313
   "010000110110000110", -- Line 1   Column 2339   Coefficient 67.38085938
   "010000110110001010", -- Line 1   Column 2340   Coefficient 67.38476563
   "010000110110001101", -- Line 1   Column 2341   Coefficient 67.38769531
   "010000110110010001", -- Line 1   Column 2342   Coefficient 67.39160156
   "010000110110010101", -- Line 1   Column 2343   Coefficient 67.39550781
   "010000110110011001", -- Line 1   Column 2344   Coefficient 67.39941406
   "010000110110011101", -- Line 1   Column 2345   Coefficient 67.40332031
   "010000110110100000", -- Line 1   Column 2346   Coefficient 67.40625000
   "010000110110100100", -- Line 1   Column 2347   Coefficient 67.41015625
   "010000110110101000", -- Line 1   Column 2348   Coefficient 67.41406250
   "010000110110101100", -- Line 1   Column 2349   Coefficient 67.41796875
   "010000110110101111", -- Line 1   Column 2350   Coefficient 67.42089844
   "010000110110110011", -- Line 1   Column 2351   Coefficient 67.42480469
   "010000110110110111", -- Line 1   Column 2352   Coefficient 67.42871094
   "010000110110111011", -- Line 1   Column 2353   Coefficient 67.43261719
   "010000110110111111", -- Line 1   Column 2354   Coefficient 67.43652344
   "010000110111000010", -- Line 1   Column 2355   Coefficient 67.43945313
   "010000110111000110", -- Line 1   Column 2356   Coefficient 67.44335938
   "010000110111001010", -- Line 1   Column 2357   Coefficient 67.44726563
   "010000110111001110", -- Line 1   Column 2358   Coefficient 67.45117188
   "010000110111010001", -- Line 1   Column 2359   Coefficient 67.45410156
   "010000110111010101", -- Line 1   Column 2360   Coefficient 67.45800781
   "010000110111011001", -- Line 1   Column 2361   Coefficient 67.46191406
   "010000110111011101", -- Line 1   Column 2362   Coefficient 67.46582031
   "010000110111100001", -- Line 1   Column 2363   Coefficient 67.46972656
   "010000110111100100", -- Line 1   Column 2364   Coefficient 67.47265625
   "010000110111101000", -- Line 1   Column 2365   Coefficient 67.47656250
   "010000110111101100", -- Line 1   Column 2366   Coefficient 67.48046875
   "010000110111110000", -- Line 1   Column 2367   Coefficient 67.48437500
   "010000110111110011", -- Line 1   Column 2368   Coefficient 67.48730469
   "010000110111110111", -- Line 1   Column 2369   Coefficient 67.49121094
   "010000110111111011", -- Line 1   Column 2370   Coefficient 67.49511719
   "010000110111111111", -- Line 1   Column 2371   Coefficient 67.49902344
   "010000111000000010", -- Line 1   Column 2372   Coefficient 67.50195313
   "010000111000000110", -- Line 1   Column 2373   Coefficient 67.50585938
   "010000111000001010", -- Line 1   Column 2374   Coefficient 67.50976563
   "010000111000001110", -- Line 1   Column 2375   Coefficient 67.51367188
   "010000111000010001", -- Line 1   Column 2376   Coefficient 67.51660156
   "010000111000010101", -- Line 1   Column 2377   Coefficient 67.52050781
   "010000111000011001", -- Line 1   Column 2378   Coefficient 67.52441406
   "010000111000011101", -- Line 1   Column 2379   Coefficient 67.52832031
   "010000111000100000", -- Line 1   Column 2380   Coefficient 67.53125000
   "010000111000100100", -- Line 1   Column 2381   Coefficient 67.53515625
   "010000111000101000", -- Line 1   Column 2382   Coefficient 67.53906250
   "010000111000101100", -- Line 1   Column 2383   Coefficient 67.54296875
   "010000111000101111", -- Line 1   Column 2384   Coefficient 67.54589844
   "010000111000110011", -- Line 1   Column 2385   Coefficient 67.54980469
   "010000111000110111", -- Line 1   Column 2386   Coefficient 67.55371094
   "010000111000111010", -- Line 1   Column 2387   Coefficient 67.55664063
   "010000111000111110", -- Line 1   Column 2388   Coefficient 67.56054688
   "010000111001000010", -- Line 1   Column 2389   Coefficient 67.56445313
   "010000111001000110", -- Line 1   Column 2390   Coefficient 67.56835938
   "010000111001001001", -- Line 1   Column 2391   Coefficient 67.57128906
   "010000111001001101", -- Line 1   Column 2392   Coefficient 67.57519531
   "010000111001010001", -- Line 1   Column 2393   Coefficient 67.57910156
   "010000111001010100", -- Line 1   Column 2394   Coefficient 67.58203125
   "010000111001011000", -- Line 1   Column 2395   Coefficient 67.58593750
   "010000111001011100", -- Line 1   Column 2396   Coefficient 67.58984375
   "010000111001100000", -- Line 1   Column 2397   Coefficient 67.59375000
   "010000111001100011", -- Line 1   Column 2398   Coefficient 67.59667969
   "010000111001100111", -- Line 1   Column 2399   Coefficient 67.60058594
   "010000111001101011", -- Line 1   Column 2400   Coefficient 67.60449219
   "010000111001101110", -- Line 1   Column 2401   Coefficient 67.60742188
   "010000111001110010", -- Line 1   Column 2402   Coefficient 67.61132813
   "010000111001110110", -- Line 1   Column 2403   Coefficient 67.61523438
   "010000111001111010", -- Line 1   Column 2404   Coefficient 67.61914063
   "010000111001111101", -- Line 1   Column 2405   Coefficient 67.62207031
   "010000111010000001", -- Line 1   Column 2406   Coefficient 67.62597656
   "010000111010000101", -- Line 1   Column 2407   Coefficient 67.62988281
   "010000111010001000", -- Line 1   Column 2408   Coefficient 67.63281250
   "010000111010001100", -- Line 1   Column 2409   Coefficient 67.63671875
   "010000111010010000", -- Line 1   Column 2410   Coefficient 67.64062500
   "010000111010010011", -- Line 1   Column 2411   Coefficient 67.64355469
   "010000111010010111", -- Line 1   Column 2412   Coefficient 67.64746094
   "010000111010011011", -- Line 1   Column 2413   Coefficient 67.65136719
   "010000111010011110", -- Line 1   Column 2414   Coefficient 67.65429688
   "010000111010100010", -- Line 1   Column 2415   Coefficient 67.65820313
   "010000111010100110", -- Line 1   Column 2416   Coefficient 67.66210938
   "010000111010101010", -- Line 1   Column 2417   Coefficient 67.66601563
   "010000111010101101", -- Line 1   Column 2418   Coefficient 67.66894531
   "010000111010110001", -- Line 1   Column 2419   Coefficient 67.67285156
   "010000111010110101", -- Line 1   Column 2420   Coefficient 67.67675781
   "010000111010111000", -- Line 1   Column 2421   Coefficient 67.67968750
   "010000111010111100", -- Line 1   Column 2422   Coefficient 67.68359375
   "010000111011000000", -- Line 1   Column 2423   Coefficient 67.68750000
   "010000111011000011", -- Line 1   Column 2424   Coefficient 67.69042969
   "010000111011000111", -- Line 1   Column 2425   Coefficient 67.69433594
   "010000111011001011", -- Line 1   Column 2426   Coefficient 67.69824219
   "010000111011001110", -- Line 1   Column 2427   Coefficient 67.70117188
   "010000111011010010", -- Line 1   Column 2428   Coefficient 67.70507813
   "010000111011010110", -- Line 1   Column 2429   Coefficient 67.70898438
   "010000111011011001", -- Line 1   Column 2430   Coefficient 67.71191406
   "010000111011011101", -- Line 1   Column 2431   Coefficient 67.71582031
   "010000111011100001", -- Line 1   Column 2432   Coefficient 67.71972656
   "010000111011100100", -- Line 1   Column 2433   Coefficient 67.72265625
   "010000111011101000", -- Line 1   Column 2434   Coefficient 67.72656250
   "010000111011101011", -- Line 1   Column 2435   Coefficient 67.72949219
   "010000111011101111", -- Line 1   Column 2436   Coefficient 67.73339844
   "010000111011110011", -- Line 1   Column 2437   Coefficient 67.73730469
   "010000111011110110", -- Line 1   Column 2438   Coefficient 67.74023438
   "010000111011111010", -- Line 1   Column 2439   Coefficient 67.74414063
   "010000111011111110", -- Line 1   Column 2440   Coefficient 67.74804688
   "010000111100000001", -- Line 1   Column 2441   Coefficient 67.75097656
   "010000111100000101", -- Line 1   Column 2442   Coefficient 67.75488281
   "010000111100001001", -- Line 1   Column 2443   Coefficient 67.75878906
   "010000111100001100", -- Line 1   Column 2444   Coefficient 67.76171875
   "010000111100010000", -- Line 1   Column 2445   Coefficient 67.76562500
   "010000111100010100", -- Line 1   Column 2446   Coefficient 67.76953125
   "010000111100010111", -- Line 1   Column 2447   Coefficient 67.77246094
   "010000111100011011", -- Line 1   Column 2448   Coefficient 67.77636719
   "010000111100011110", -- Line 1   Column 2449   Coefficient 67.77929688
   "010000111100100010", -- Line 1   Column 2450   Coefficient 67.78320313
   "010000111100100110", -- Line 1   Column 2451   Coefficient 67.78710938
   "010000111100101001", -- Line 1   Column 2452   Coefficient 67.79003906
   "010000111100101101", -- Line 1   Column 2453   Coefficient 67.79394531
   "010000111100110001", -- Line 1   Column 2454   Coefficient 67.79785156
   "010000111100110100", -- Line 1   Column 2455   Coefficient 67.80078125
   "010000111100111000", -- Line 1   Column 2456   Coefficient 67.80468750
   "010000111100111011", -- Line 1   Column 2457   Coefficient 67.80761719
   "010000111100111111", -- Line 1   Column 2458   Coefficient 67.81152344
   "010000111101000011", -- Line 1   Column 2459   Coefficient 67.81542969
   "010000111101000110", -- Line 1   Column 2460   Coefficient 67.81835938
   "010000111101001010", -- Line 1   Column 2461   Coefficient 67.82226563
   "010000111101001110", -- Line 1   Column 2462   Coefficient 67.82617188
   "010000111101010001", -- Line 1   Column 2463   Coefficient 67.82910156
   "010000111101010101", -- Line 1   Column 2464   Coefficient 67.83300781
   "010000111101011000", -- Line 1   Column 2465   Coefficient 67.83593750
   "010000111101011100", -- Line 1   Column 2466   Coefficient 67.83984375
   "010000111101100000", -- Line 1   Column 2467   Coefficient 67.84375000
   "010000111101100011", -- Line 1   Column 2468   Coefficient 67.84667969
   "010000111101100111", -- Line 1   Column 2469   Coefficient 67.85058594
   "010000111101101010", -- Line 1   Column 2470   Coefficient 67.85351563
   "010000111101101110", -- Line 1   Column 2471   Coefficient 67.85742188
   "010000111101110010", -- Line 1   Column 2472   Coefficient 67.86132813
   "010000111101110101", -- Line 1   Column 2473   Coefficient 67.86425781
   "010000111101111001", -- Line 1   Column 2474   Coefficient 67.86816406
   "010000111101111100", -- Line 1   Column 2475   Coefficient 67.87109375
   "010000111110000000", -- Line 1   Column 2476   Coefficient 67.87500000
   "010000111110000100", -- Line 1   Column 2477   Coefficient 67.87890625
   "010000111110000111", -- Line 1   Column 2478   Coefficient 67.88183594
   "010000111110001011", -- Line 1   Column 2479   Coefficient 67.88574219
   "010000111110001110", -- Line 1   Column 2480   Coefficient 67.88867188
   "010000111110010010", -- Line 1   Column 2481   Coefficient 67.89257813
   "010000111110010110", -- Line 1   Column 2482   Coefficient 67.89648438
   "010000111110011001", -- Line 1   Column 2483   Coefficient 67.89941406
   "010000111110011101", -- Line 1   Column 2484   Coefficient 67.90332031
   "010000111110100000", -- Line 1   Column 2485   Coefficient 67.90625000
   "010000111110100100", -- Line 1   Column 2486   Coefficient 67.91015625
   "010000111110100111", -- Line 1   Column 2487   Coefficient 67.91308594
   "010000111110101011", -- Line 1   Column 2488   Coefficient 67.91699219
   "010000111110101111", -- Line 1   Column 2489   Coefficient 67.92089844
   "010000111110110010", -- Line 1   Column 2490   Coefficient 67.92382813
   "010000111110110110", -- Line 1   Column 2491   Coefficient 67.92773438
   "010000111110111001", -- Line 1   Column 2492   Coefficient 67.93066406
   "010000111110111101", -- Line 1   Column 2493   Coefficient 67.93457031
   "010000111111000000", -- Line 1   Column 2494   Coefficient 67.93750000
   "010000111111000100", -- Line 1   Column 2495   Coefficient 67.94140625
   "010000111111001000", -- Line 1   Column 2496   Coefficient 67.94531250
   "010000111111001011", -- Line 1   Column 2497   Coefficient 67.94824219
   "010000111111001111", -- Line 1   Column 2498   Coefficient 67.95214844
   "010000111111010010", -- Line 1   Column 2499   Coefficient 67.95507813
   "010000111111010110", -- Line 1   Column 2500   Coefficient 67.95898438
   "010000111111011001", -- Line 1   Column 2501   Coefficient 67.96191406
   "010000111111011101", -- Line 1   Column 2502   Coefficient 67.96582031
   "010000111111100000", -- Line 1   Column 2503   Coefficient 67.96875000
   "010000111111100100", -- Line 1   Column 2504   Coefficient 67.97265625
   "010000111111101000", -- Line 1   Column 2505   Coefficient 67.97656250
   "010000111111101011", -- Line 1   Column 2506   Coefficient 67.97949219
   "010000111111101111", -- Line 1   Column 2507   Coefficient 67.98339844
   "010000111111110010", -- Line 1   Column 2508   Coefficient 67.98632813
   "010000111111110110", -- Line 1   Column 2509   Coefficient 67.99023438
   "010000111111111001", -- Line 1   Column 2510   Coefficient 67.99316406
   "010000111111111101", -- Line 1   Column 2511   Coefficient 67.99707031
   "010001000000000000", -- Line 1   Column 2512   Coefficient 68.00000000
   "010001000000000100", -- Line 1   Column 2513   Coefficient 68.00390625
   "010001000000000111", -- Line 1   Column 2514   Coefficient 68.00683594
   "010001000000001011", -- Line 1   Column 2515   Coefficient 68.01074219
   "010001000000001111", -- Line 1   Column 2516   Coefficient 68.01464844
   "010001000000010010", -- Line 1   Column 2517   Coefficient 68.01757813
   "010001000000010110", -- Line 1   Column 2518   Coefficient 68.02148438
   "010001000000011001", -- Line 1   Column 2519   Coefficient 68.02441406
   "010001000000011101", -- Line 1   Column 2520   Coefficient 68.02832031
   "010001000000100000", -- Line 1   Column 2521   Coefficient 68.03125000
   "010001000000100100", -- Line 1   Column 2522   Coefficient 68.03515625
   "010001000000100111", -- Line 1   Column 2523   Coefficient 68.03808594
   "010001000000101011", -- Line 1   Column 2524   Coefficient 68.04199219
   "010001000000101110", -- Line 1   Column 2525   Coefficient 68.04492188
   "010001000000110010", -- Line 1   Column 2526   Coefficient 68.04882813
   "010001000000110101", -- Line 1   Column 2527   Coefficient 68.05175781
   "010001000000111001", -- Line 1   Column 2528   Coefficient 68.05566406
   "010001000000111100", -- Line 1   Column 2529   Coefficient 68.05859375
   "010001000001000000", -- Line 1   Column 2530   Coefficient 68.06250000
   "010001000001000011", -- Line 1   Column 2531   Coefficient 68.06542969
   "010001000001000111", -- Line 1   Column 2532   Coefficient 68.06933594
   "010001000001001010", -- Line 1   Column 2533   Coefficient 68.07226563
   "010001000001001110", -- Line 1   Column 2534   Coefficient 68.07617188
   "010001000001010001", -- Line 1   Column 2535   Coefficient 68.07910156
   "010001000001010101", -- Line 1   Column 2536   Coefficient 68.08300781
   "010001000001011000", -- Line 1   Column 2537   Coefficient 68.08593750
   "010001000001011100", -- Line 1   Column 2538   Coefficient 68.08984375
   "010001000001011111", -- Line 1   Column 2539   Coefficient 68.09277344
   "010001000001100011", -- Line 1   Column 2540   Coefficient 68.09667969
   "010001000001100110", -- Line 1   Column 2541   Coefficient 68.09960938
   "010001000001101010", -- Line 1   Column 2542   Coefficient 68.10351563
   "010001000001101101", -- Line 1   Column 2543   Coefficient 68.10644531
   "010001000001110001", -- Line 1   Column 2544   Coefficient 68.11035156
   "010001000001110100", -- Line 1   Column 2545   Coefficient 68.11328125
   "010001000001111000", -- Line 1   Column 2546   Coefficient 68.11718750
   "010001000001111011", -- Line 1   Column 2547   Coefficient 68.12011719
   "010001000001111111", -- Line 1   Column 2548   Coefficient 68.12402344
   "010001000010000010", -- Line 1   Column 2549   Coefficient 68.12695313
   "010001000010000110", -- Line 1   Column 2550   Coefficient 68.13085938
   "010001000010001001", -- Line 1   Column 2551   Coefficient 68.13378906
   "010001000010001101", -- Line 1   Column 2552   Coefficient 68.13769531
   "010001000010010000", -- Line 1   Column 2553   Coefficient 68.14062500
   "010001000010010100", -- Line 1   Column 2554   Coefficient 68.14453125
   "010001000010010111", -- Line 1   Column 2555   Coefficient 68.14746094
   "010001000010011011", -- Line 1   Column 2556   Coefficient 68.15136719
   "010001000010011110", -- Line 1   Column 2557   Coefficient 68.15429688
   "010001000010100010", -- Line 1   Column 2558   Coefficient 68.15820313
   "010001000010100101", -- Line 1   Column 2559   Coefficient 68.16113281
   "010001000010101001", -- Line 1   Column 2560   Coefficient 68.16503906
   "010001000010101100", -- Line 1   Column 2561   Coefficient 68.16796875
   "010001000010110000", -- Line 1   Column 2562   Coefficient 68.17187500
   "010001000010110011", -- Line 1   Column 2563   Coefficient 68.17480469
   "010001000010110111", -- Line 1   Column 2564   Coefficient 68.17871094
   "010001000010111010", -- Line 1   Column 2565   Coefficient 68.18164063
   "010001000010111110", -- Line 1   Column 2566   Coefficient 68.18554688
   "010001000011000001", -- Line 1   Column 2567   Coefficient 68.18847656
   "010001000011000101", -- Line 1   Column 2568   Coefficient 68.19238281
   "010001000011001000", -- Line 1   Column 2569   Coefficient 68.19531250
   "010001000011001011", -- Line 1   Column 2570   Coefficient 68.19824219
   "010001000011001111", -- Line 1   Column 2571   Coefficient 68.20214844
   "010001000011010010", -- Line 1   Column 2572   Coefficient 68.20507813
   "010001000011010110", -- Line 1   Column 2573   Coefficient 68.20898438
   "010001000011011001", -- Line 1   Column 2574   Coefficient 68.21191406
   "010001000011011101", -- Line 1   Column 2575   Coefficient 68.21582031
   "010001000011100000", -- Line 1   Column 2576   Coefficient 68.21875000
   "010001000011100100", -- Line 1   Column 2577   Coefficient 68.22265625
   "010001000011100111", -- Line 1   Column 2578   Coefficient 68.22558594
   "010001000011101011", -- Line 1   Column 2579   Coefficient 68.22949219
   "010001000011101110", -- Line 1   Column 2580   Coefficient 68.23242188
   "010001000011110001", -- Line 1   Column 2581   Coefficient 68.23535156
   "010001000011110101", -- Line 1   Column 2582   Coefficient 68.23925781
   "010001000011111000", -- Line 1   Column 2583   Coefficient 68.24218750
   "010001000011111100", -- Line 1   Column 2584   Coefficient 68.24609375
   "010001000011111111", -- Line 1   Column 2585   Coefficient 68.24902344
   "010001000100000011", -- Line 1   Column 2586   Coefficient 68.25292969
   "010001000100000110", -- Line 1   Column 2587   Coefficient 68.25585938
   "010001000100001010", -- Line 1   Column 2588   Coefficient 68.25976563
   "010001000100001101", -- Line 1   Column 2589   Coefficient 68.26269531
   "010001000100010000", -- Line 1   Column 2590   Coefficient 68.26562500
   "010001000100010100", -- Line 1   Column 2591   Coefficient 68.26953125
   "010001000100010111", -- Line 1   Column 2592   Coefficient 68.27246094
   "010001000100011011", -- Line 1   Column 2593   Coefficient 68.27636719
   "010001000100011110", -- Line 1   Column 2594   Coefficient 68.27929688
   "010001000100100010", -- Line 1   Column 2595   Coefficient 68.28320313
   "010001000100100101", -- Line 1   Column 2596   Coefficient 68.28613281
   "010001000100101000", -- Line 1   Column 2597   Coefficient 68.28906250
   "010001000100101100", -- Line 1   Column 2598   Coefficient 68.29296875
   "010001000100101111", -- Line 1   Column 2599   Coefficient 68.29589844
   "010001000100110011", -- Line 1   Column 2600   Coefficient 68.29980469
   "010001000100110110", -- Line 1   Column 2601   Coefficient 68.30273438
   "010001000100111001", -- Line 1   Column 2602   Coefficient 68.30566406
   "010001000100111101", -- Line 1   Column 2603   Coefficient 68.30957031
   "010001000101000000", -- Line 1   Column 2604   Coefficient 68.31250000
   "010001000101000100", -- Line 1   Column 2605   Coefficient 68.31640625
   "010001000101000111", -- Line 1   Column 2606   Coefficient 68.31933594
   "010001000101001011", -- Line 1   Column 2607   Coefficient 68.32324219
   "010001000101001110", -- Line 1   Column 2608   Coefficient 68.32617188
   "010001000101010001", -- Line 1   Column 2609   Coefficient 68.32910156
   "010001000101010101", -- Line 1   Column 2610   Coefficient 68.33300781
   "010001000101011000", -- Line 1   Column 2611   Coefficient 68.33593750
   "010001000101011100", -- Line 1   Column 2612   Coefficient 68.33984375
   "010001000101011111", -- Line 1   Column 2613   Coefficient 68.34277344
   "010001000101100010", -- Line 1   Column 2614   Coefficient 68.34570313
   "010001000101100110", -- Line 1   Column 2615   Coefficient 68.34960938
   "010001000101101001", -- Line 1   Column 2616   Coefficient 68.35253906
   "010001000101101101", -- Line 1   Column 2617   Coefficient 68.35644531
   "010001000101110000", -- Line 1   Column 2618   Coefficient 68.35937500
   "010001000101110011", -- Line 1   Column 2619   Coefficient 68.36230469
   "010001000101110111", -- Line 1   Column 2620   Coefficient 68.36621094
   "010001000101111010", -- Line 1   Column 2621   Coefficient 68.36914063
   "010001000101111110", -- Line 1   Column 2622   Coefficient 68.37304688
   "010001000110000001", -- Line 1   Column 2623   Coefficient 68.37597656
   "010001000110000100", -- Line 1   Column 2624   Coefficient 68.37890625
   "010001000110001000", -- Line 1   Column 2625   Coefficient 68.38281250
   "010001000110001011", -- Line 1   Column 2626   Coefficient 68.38574219
   "010001000110001111", -- Line 1   Column 2627   Coefficient 68.38964844
   "010001000110010010", -- Line 1   Column 2628   Coefficient 68.39257813
   "010001000110010101", -- Line 1   Column 2629   Coefficient 68.39550781
   "010001000110011001", -- Line 1   Column 2630   Coefficient 68.39941406
   "010001000110011100", -- Line 1   Column 2631   Coefficient 68.40234375
   "010001000110011111", -- Line 1   Column 2632   Coefficient 68.40527344
   "010001000110100011", -- Line 1   Column 2633   Coefficient 68.40917969
   "010001000110100110", -- Line 1   Column 2634   Coefficient 68.41210938
   "010001000110101010", -- Line 1   Column 2635   Coefficient 68.41601563
   "010001000110101101", -- Line 1   Column 2636   Coefficient 68.41894531
   "010001000110110000", -- Line 1   Column 2637   Coefficient 68.42187500
   "010001000110110100", -- Line 1   Column 2638   Coefficient 68.42578125
   "010001000110110111", -- Line 1   Column 2639   Coefficient 68.42871094
   "010001000110111010", -- Line 1   Column 2640   Coefficient 68.43164063
   "010001000110111110", -- Line 1   Column 2641   Coefficient 68.43554688
   "010001000111000001", -- Line 1   Column 2642   Coefficient 68.43847656
   "010001000111000101", -- Line 1   Column 2643   Coefficient 68.44238281
   "010001000111001000", -- Line 1   Column 2644   Coefficient 68.44531250
   "010001000111001011", -- Line 1   Column 2645   Coefficient 68.44824219
   "010001000111001111", -- Line 1   Column 2646   Coefficient 68.45214844
   "010001000111010010", -- Line 1   Column 2647   Coefficient 68.45507813
   "010001000111010101", -- Line 1   Column 2648   Coefficient 68.45800781
   "010001000111011001", -- Line 1   Column 2649   Coefficient 68.46191406
   "010001000111011100", -- Line 1   Column 2650   Coefficient 68.46484375
   "010001000111011111", -- Line 1   Column 2651   Coefficient 68.46777344
   "010001000111100011", -- Line 1   Column 2652   Coefficient 68.47167969
   "010001000111100110", -- Line 1   Column 2653   Coefficient 68.47460938
   "010001000111101001", -- Line 1   Column 2654   Coefficient 68.47753906
   "010001000111101101", -- Line 1   Column 2655   Coefficient 68.48144531
   "010001000111110000", -- Line 1   Column 2656   Coefficient 68.48437500
   "010001000111110100", -- Line 1   Column 2657   Coefficient 68.48828125
   "010001000111110111", -- Line 1   Column 2658   Coefficient 68.49121094
   "010001000111111010", -- Line 1   Column 2659   Coefficient 68.49414063
   "010001000111111110", -- Line 1   Column 2660   Coefficient 68.49804688
   "010001001000000001", -- Line 1   Column 2661   Coefficient 68.50097656
   "010001001000000100", -- Line 1   Column 2662   Coefficient 68.50390625
   "010001001000001000", -- Line 1   Column 2663   Coefficient 68.50781250
   "010001001000001011", -- Line 1   Column 2664   Coefficient 68.51074219
   "010001001000001110", -- Line 1   Column 2665   Coefficient 68.51367188
   "010001001000010010", -- Line 1   Column 2666   Coefficient 68.51757813
   "010001001000010101", -- Line 1   Column 2667   Coefficient 68.52050781
   "010001001000011000", -- Line 1   Column 2668   Coefficient 68.52343750
   "010001001000011100", -- Line 1   Column 2669   Coefficient 68.52734375
   "010001001000011111", -- Line 1   Column 2670   Coefficient 68.53027344
   "010001001000100010", -- Line 1   Column 2671   Coefficient 68.53320313
   "010001001000100110", -- Line 1   Column 2672   Coefficient 68.53710938
   "010001001000101001", -- Line 1   Column 2673   Coefficient 68.54003906
   "010001001000101100", -- Line 1   Column 2674   Coefficient 68.54296875
   "010001001000110000", -- Line 1   Column 2675   Coefficient 68.54687500
   "010001001000110011", -- Line 1   Column 2676   Coefficient 68.54980469
   "010001001000110110", -- Line 1   Column 2677   Coefficient 68.55273438
   "010001001000111010", -- Line 1   Column 2678   Coefficient 68.55664063
   "010001001000111101", -- Line 1   Column 2679   Coefficient 68.55957031
   "010001001001000000", -- Line 1   Column 2680   Coefficient 68.56250000
   "010001001001000100", -- Line 1   Column 2681   Coefficient 68.56640625
   "010001001001000111", -- Line 1   Column 2682   Coefficient 68.56933594
   "010001001001001010", -- Line 1   Column 2683   Coefficient 68.57226563
   "010001001001001101", -- Line 1   Column 2684   Coefficient 68.57519531
   "010001001001010001", -- Line 1   Column 2685   Coefficient 68.57910156
   "010001001001010100", -- Line 1   Column 2686   Coefficient 68.58203125
   "010001001001010111", -- Line 1   Column 2687   Coefficient 68.58496094
   "010001001001011011", -- Line 1   Column 2688   Coefficient 68.58886719
   "010001001001011110", -- Line 1   Column 2689   Coefficient 68.59179688
   "010001001001100001", -- Line 1   Column 2690   Coefficient 68.59472656
   "010001001001100101", -- Line 1   Column 2691   Coefficient 68.59863281
   "010001001001101000", -- Line 1   Column 2692   Coefficient 68.60156250
   "010001001001101011", -- Line 1   Column 2693   Coefficient 68.60449219
   "010001001001101111", -- Line 1   Column 2694   Coefficient 68.60839844
   "010001001001110010", -- Line 1   Column 2695   Coefficient 68.61132813
   "010001001001110101", -- Line 1   Column 2696   Coefficient 68.61425781
   "010001001001111000", -- Line 1   Column 2697   Coefficient 68.61718750
   "010001001001111100", -- Line 1   Column 2698   Coefficient 68.62109375
   "010001001001111111", -- Line 1   Column 2699   Coefficient 68.62402344
   "010001001010000010", -- Line 1   Column 2700   Coefficient 68.62695313
   "010001001010000110", -- Line 1   Column 2701   Coefficient 68.63085938
   "010001001010001001", -- Line 1   Column 2702   Coefficient 68.63378906
   "010001001010001100", -- Line 1   Column 2703   Coefficient 68.63671875
   "010001001010001111", -- Line 1   Column 2704   Coefficient 68.63964844
   "010001001010010011", -- Line 1   Column 2705   Coefficient 68.64355469
   "010001001010010110", -- Line 1   Column 2706   Coefficient 68.64648438
   "010001001010011001", -- Line 1   Column 2707   Coefficient 68.64941406
   "010001001010011101", -- Line 1   Column 2708   Coefficient 68.65332031
   "010001001010100000", -- Line 1   Column 2709   Coefficient 68.65625000
   "010001001010100011", -- Line 1   Column 2710   Coefficient 68.65917969
   "010001001010100110", -- Line 1   Column 2711   Coefficient 68.66210938
   "010001001010101010", -- Line 1   Column 2712   Coefficient 68.66601563
   "010001001010101101", -- Line 1   Column 2713   Coefficient 68.66894531
   "010001001010110000", -- Line 1   Column 2714   Coefficient 68.67187500
   "010001001010110100", -- Line 1   Column 2715   Coefficient 68.67578125
   "010001001010110111", -- Line 1   Column 2716   Coefficient 68.67871094
   "010001001010111010", -- Line 1   Column 2717   Coefficient 68.68164063
   "010001001010111101", -- Line 1   Column 2718   Coefficient 68.68457031
   "010001001011000001", -- Line 1   Column 2719   Coefficient 68.68847656
   "010001001011000100", -- Line 1   Column 2720   Coefficient 68.69140625
   "010001001011000111", -- Line 1   Column 2721   Coefficient 68.69433594
   "010001001011001011", -- Line 1   Column 2722   Coefficient 68.69824219
   "010001001011001110", -- Line 1   Column 2723   Coefficient 68.70117188
   "010001001011010001", -- Line 1   Column 2724   Coefficient 68.70410156
   "010001001011010100", -- Line 1   Column 2725   Coefficient 68.70703125
   "010001001011011000", -- Line 1   Column 2726   Coefficient 68.71093750
   "010001001011011011", -- Line 1   Column 2727   Coefficient 68.71386719
   "010001001011011110", -- Line 1   Column 2728   Coefficient 68.71679688
   "010001001011100001", -- Line 1   Column 2729   Coefficient 68.71972656
   "010001001011100101", -- Line 1   Column 2730   Coefficient 68.72363281
   "010001001011101000", -- Line 1   Column 2731   Coefficient 68.72656250
   "010001001011101011", -- Line 1   Column 2732   Coefficient 68.72949219
   "010001001011101110", -- Line 1   Column 2733   Coefficient 68.73242188
   "010001001011110010", -- Line 1   Column 2734   Coefficient 68.73632813
   "010001001011110101", -- Line 1   Column 2735   Coefficient 68.73925781
   "010001001011111000", -- Line 1   Column 2736   Coefficient 68.74218750
   "010001001011111011", -- Line 1   Column 2737   Coefficient 68.74511719
   "010001001011111111", -- Line 1   Column 2738   Coefficient 68.74902344
   "010001001100000010", -- Line 1   Column 2739   Coefficient 68.75195313
   "010001001100000101", -- Line 1   Column 2740   Coefficient 68.75488281
   "010001001100001000", -- Line 1   Column 2741   Coefficient 68.75781250
   "010001001100001100", -- Line 1   Column 2742   Coefficient 68.76171875
   "010001001100001111", -- Line 1   Column 2743   Coefficient 68.76464844
   "010001001100010010", -- Line 1   Column 2744   Coefficient 68.76757813
   "010001001100010101", -- Line 1   Column 2745   Coefficient 68.77050781
   "010001001100011001", -- Line 1   Column 2746   Coefficient 68.77441406
   "010001001100011100", -- Line 1   Column 2747   Coefficient 68.77734375
   "010001001100011111", -- Line 1   Column 2748   Coefficient 68.78027344
   "010001001100100010", -- Line 1   Column 2749   Coefficient 68.78320313
   "010001001100100110", -- Line 1   Column 2750   Coefficient 68.78710938
   "010001001100101001", -- Line 1   Column 2751   Coefficient 68.79003906
   "010001001100101100", -- Line 1   Column 2752   Coefficient 68.79296875
   "010001001100101111", -- Line 1   Column 2753   Coefficient 68.79589844
   "010001001100110010", -- Line 1   Column 2754   Coefficient 68.79882813
   "010001001100110110", -- Line 1   Column 2755   Coefficient 68.80273438
   "010001001100111001", -- Line 1   Column 2756   Coefficient 68.80566406
   "010001001100111100", -- Line 1   Column 2757   Coefficient 68.80859375
   "010001001100111111", -- Line 1   Column 2758   Coefficient 68.81152344
   "010001001101000011", -- Line 1   Column 2759   Coefficient 68.81542969
   "010001001101000110", -- Line 1   Column 2760   Coefficient 68.81835938
   "010001001101001001", -- Line 1   Column 2761   Coefficient 68.82128906
   "010001001101001100", -- Line 1   Column 2762   Coefficient 68.82421875
   "010001001101001111", -- Line 1   Column 2763   Coefficient 68.82714844
   "010001001101010011", -- Line 1   Column 2764   Coefficient 68.83105469
   "010001001101010110", -- Line 1   Column 2765   Coefficient 68.83398438
   "010001001101011001", -- Line 1   Column 2766   Coefficient 68.83691406
   "010001001101011100", -- Line 1   Column 2767   Coefficient 68.83984375
   "010001001101100000", -- Line 1   Column 2768   Coefficient 68.84375000
   "010001001101100011", -- Line 1   Column 2769   Coefficient 68.84667969
   "010001001101100110", -- Line 1   Column 2770   Coefficient 68.84960938
   "010001001101101001", -- Line 1   Column 2771   Coefficient 68.85253906
   "010001001101101100", -- Line 1   Column 2772   Coefficient 68.85546875
   "010001001101110000", -- Line 1   Column 2773   Coefficient 68.85937500
   "010001001101110011", -- Line 1   Column 2774   Coefficient 68.86230469
   "010001001101110110", -- Line 1   Column 2775   Coefficient 68.86523438
   "010001001101111001", -- Line 1   Column 2776   Coefficient 68.86816406
   "010001001101111100", -- Line 1   Column 2777   Coefficient 68.87109375
   "010001001110000000", -- Line 1   Column 2778   Coefficient 68.87500000
   "010001001110000011", -- Line 1   Column 2779   Coefficient 68.87792969
   "010001001110000110", -- Line 1   Column 2780   Coefficient 68.88085938
   "010001001110001001", -- Line 1   Column 2781   Coefficient 68.88378906
   "010001001110001100", -- Line 1   Column 2782   Coefficient 68.88671875
   "010001001110010000", -- Line 1   Column 2783   Coefficient 68.89062500
   "010001001110010011", -- Line 1   Column 2784   Coefficient 68.89355469
   "010001001110010110", -- Line 1   Column 2785   Coefficient 68.89648438
   "010001001110011001", -- Line 1   Column 2786   Coefficient 68.89941406
   "010001001110011100", -- Line 1   Column 2787   Coefficient 68.90234375
   "010001001110100000", -- Line 1   Column 2788   Coefficient 68.90625000
   "010001001110100011", -- Line 1   Column 2789   Coefficient 68.90917969
   "010001001110100110", -- Line 1   Column 2790   Coefficient 68.91210938
   "010001001110101001", -- Line 1   Column 2791   Coefficient 68.91503906
   "010001001110101100", -- Line 1   Column 2792   Coefficient 68.91796875
   "010001001110110000", -- Line 1   Column 2793   Coefficient 68.92187500
   "010001001110110011", -- Line 1   Column 2794   Coefficient 68.92480469
   "010001001110110110", -- Line 1   Column 2795   Coefficient 68.92773438
   "010001001110111001", -- Line 1   Column 2796   Coefficient 68.93066406
   "010001001110111100", -- Line 1   Column 2797   Coefficient 68.93359375
   "010001001110111111", -- Line 1   Column 2798   Coefficient 68.93652344
   "010001001111000011", -- Line 1   Column 2799   Coefficient 68.94042969
   "010001001111000110", -- Line 1   Column 2800   Coefficient 68.94335938
   "010001001111001001", -- Line 1   Column 2801   Coefficient 68.94628906
   "010001001111001100", -- Line 1   Column 2802   Coefficient 68.94921875
   "010001001111001111", -- Line 1   Column 2803   Coefficient 68.95214844
   "010001001111010010", -- Line 1   Column 2804   Coefficient 68.95507813
   "010001001111010110", -- Line 1   Column 2805   Coefficient 68.95898438
   "010001001111011001", -- Line 1   Column 2806   Coefficient 68.96191406
   "010001001111011100", -- Line 1   Column 2807   Coefficient 68.96484375
   "010001001111011111", -- Line 1   Column 2808   Coefficient 68.96777344
   "010001001111100010", -- Line 1   Column 2809   Coefficient 68.97070313
   "010001001111100110", -- Line 1   Column 2810   Coefficient 68.97460938
   "010001001111101001", -- Line 1   Column 2811   Coefficient 68.97753906
   "010001001111101100", -- Line 1   Column 2812   Coefficient 68.98046875
   "010001001111101111", -- Line 1   Column 2813   Coefficient 68.98339844
   "010001001111110010", -- Line 1   Column 2814   Coefficient 68.98632813
   "010001001111110101", -- Line 1   Column 2815   Coefficient 68.98925781
   "010001001111111000", -- Line 1   Column 2816   Coefficient 68.99218750
   "010001001111111100", -- Line 1   Column 2817   Coefficient 68.99609375
   "010001001111111111", -- Line 1   Column 2818   Coefficient 68.99902344
   "010001010000000010", -- Line 1   Column 2819   Coefficient 69.00195313
   "010001010000000101", -- Line 1   Column 2820   Coefficient 69.00488281
   "010001010000001000", -- Line 1   Column 2821   Coefficient 69.00781250
   "010001010000001011", -- Line 1   Column 2822   Coefficient 69.01074219
   "010001010000001111", -- Line 1   Column 2823   Coefficient 69.01464844
   "010001010000010010", -- Line 1   Column 2824   Coefficient 69.01757813
   "010001010000010101", -- Line 1   Column 2825   Coefficient 69.02050781
   "010001010000011000", -- Line 1   Column 2826   Coefficient 69.02343750
   "010001010000011011", -- Line 1   Column 2827   Coefficient 69.02636719
   "010001010000011110", -- Line 1   Column 2828   Coefficient 69.02929688
   "010001010000100001", -- Line 1   Column 2829   Coefficient 69.03222656
   "010001010000100101", -- Line 1   Column 2830   Coefficient 69.03613281
   "010001010000101000", -- Line 1   Column 2831   Coefficient 69.03906250
   "010001010000101011", -- Line 1   Column 2832   Coefficient 69.04199219
   "010001010000101110", -- Line 1   Column 2833   Coefficient 69.04492188
   "010001010000110001", -- Line 1   Column 2834   Coefficient 69.04785156
   "010001010000110100", -- Line 1   Column 2835   Coefficient 69.05078125
   "010001010000110111", -- Line 1   Column 2836   Coefficient 69.05371094
   "010001010000111011", -- Line 1   Column 2837   Coefficient 69.05761719
   "010001010000111110", -- Line 1   Column 2838   Coefficient 69.06054688
   "010001010001000001", -- Line 1   Column 2839   Coefficient 69.06347656
   "010001010001000100", -- Line 1   Column 2840   Coefficient 69.06640625
   "010001010001000111", -- Line 1   Column 2841   Coefficient 69.06933594
   "010001010001001010", -- Line 1   Column 2842   Coefficient 69.07226563
   "010001010001001101", -- Line 1   Column 2843   Coefficient 69.07519531
   "010001010001010000", -- Line 1   Column 2844   Coefficient 69.07812500
   "010001010001010100", -- Line 1   Column 2845   Coefficient 69.08203125
   "010001010001010111", -- Line 1   Column 2846   Coefficient 69.08496094
   "010001010001011010", -- Line 1   Column 2847   Coefficient 69.08789063
   "010001010001011101", -- Line 1   Column 2848   Coefficient 69.09082031
   "010001010001100000", -- Line 1   Column 2849   Coefficient 69.09375000
   "010001010001100011", -- Line 1   Column 2850   Coefficient 69.09667969
   "010001010001100110", -- Line 1   Column 2851   Coefficient 69.09960938
   "010001010001101001", -- Line 1   Column 2852   Coefficient 69.10253906
   "010001010001101101", -- Line 1   Column 2853   Coefficient 69.10644531
   "010001010001110000", -- Line 1   Column 2854   Coefficient 69.10937500
   "010001010001110011", -- Line 1   Column 2855   Coefficient 69.11230469
   "010001010001110110", -- Line 1   Column 2856   Coefficient 69.11523438
   "010001010001111001", -- Line 1   Column 2857   Coefficient 69.11816406
   "010001010001111100", -- Line 1   Column 2858   Coefficient 69.12109375
   "010001010001111111", -- Line 1   Column 2859   Coefficient 69.12402344
   "010001010010000010", -- Line 1   Column 2860   Coefficient 69.12695313
   "010001010010000101", -- Line 1   Column 2861   Coefficient 69.12988281
   "010001010010001001", -- Line 1   Column 2862   Coefficient 69.13378906
   "010001010010001100", -- Line 1   Column 2863   Coefficient 69.13671875
   "010001010010001111", -- Line 1   Column 2864   Coefficient 69.13964844
   "010001010010010010", -- Line 1   Column 2865   Coefficient 69.14257813
   "010001010010010101", -- Line 1   Column 2866   Coefficient 69.14550781
   "010001010010011000", -- Line 1   Column 2867   Coefficient 69.14843750
   "010001010010011011", -- Line 1   Column 2868   Coefficient 69.15136719
   "010001010010011110", -- Line 1   Column 2869   Coefficient 69.15429688
   "010001010010100001", -- Line 1   Column 2870   Coefficient 69.15722656
   "010001010010100101", -- Line 1   Column 2871   Coefficient 69.16113281
   "010001010010101000", -- Line 1   Column 2872   Coefficient 69.16406250
   "010001010010101011", -- Line 1   Column 2873   Coefficient 69.16699219
   "010001010010101110", -- Line 1   Column 2874   Coefficient 69.16992188
   "010001010010110001", -- Line 1   Column 2875   Coefficient 69.17285156
   "010001010010110100", -- Line 1   Column 2876   Coefficient 69.17578125
   "010001010010110111", -- Line 1   Column 2877   Coefficient 69.17871094
   "010001010010111010", -- Line 1   Column 2878   Coefficient 69.18164063
   "010001010010111101", -- Line 1   Column 2879   Coefficient 69.18457031
   "010001010011000000", -- Line 1   Column 2880   Coefficient 69.18750000
   "010001010011000011", -- Line 1   Column 2881   Coefficient 69.19042969
   "010001010011000111", -- Line 1   Column 2882   Coefficient 69.19433594
   "010001010011001010", -- Line 1   Column 2883   Coefficient 69.19726563
   "010001010011001101", -- Line 1   Column 2884   Coefficient 69.20019531
   "010001010011010000", -- Line 1   Column 2885   Coefficient 69.20312500
   "010001010011010011", -- Line 1   Column 2886   Coefficient 69.20605469
   "010001010011010110", -- Line 1   Column 2887   Coefficient 69.20898438
   "010001010011011001", -- Line 1   Column 2888   Coefficient 69.21191406
   "010001010011011100", -- Line 1   Column 2889   Coefficient 69.21484375
   "010001010011011111", -- Line 1   Column 2890   Coefficient 69.21777344
   "010001010011100010", -- Line 1   Column 2891   Coefficient 69.22070313
   "010001010011100101", -- Line 1   Column 2892   Coefficient 69.22363281
   "010001010011101000", -- Line 1   Column 2893   Coefficient 69.22656250
   "010001010011101011", -- Line 1   Column 2894   Coefficient 69.22949219
   "010001010011101111", -- Line 1   Column 2895   Coefficient 69.23339844
   "010001010011110010", -- Line 1   Column 2896   Coefficient 69.23632813
   "010001010011110101", -- Line 1   Column 2897   Coefficient 69.23925781
   "010001010011111000", -- Line 1   Column 2898   Coefficient 69.24218750
   "010001010011111011", -- Line 1   Column 2899   Coefficient 69.24511719
   "010001010011111110", -- Line 1   Column 2900   Coefficient 69.24804688
   "010001010100000001", -- Line 1   Column 2901   Coefficient 69.25097656
   "010001010100000100", -- Line 1   Column 2902   Coefficient 69.25390625
   "010001010100000111", -- Line 1   Column 2903   Coefficient 69.25683594
   "010001010100001010", -- Line 1   Column 2904   Coefficient 69.25976563
   "010001010100001101", -- Line 1   Column 2905   Coefficient 69.26269531
   "010001010100010000", -- Line 1   Column 2906   Coefficient 69.26562500
   "010001010100010011", -- Line 1   Column 2907   Coefficient 69.26855469
   "010001010100010110", -- Line 1   Column 2908   Coefficient 69.27148438
   "010001010100011001", -- Line 1   Column 2909   Coefficient 69.27441406
   "010001010100011101", -- Line 1   Column 2910   Coefficient 69.27832031
   "010001010100100000", -- Line 1   Column 2911   Coefficient 69.28125000
   "010001010100100011", -- Line 1   Column 2912   Coefficient 69.28417969
   "010001010100100110", -- Line 1   Column 2913   Coefficient 69.28710938
   "010001010100101001", -- Line 1   Column 2914   Coefficient 69.29003906
   "010001010100101100", -- Line 1   Column 2915   Coefficient 69.29296875
   "010001010100101111", -- Line 1   Column 2916   Coefficient 69.29589844
   "010001010100110010", -- Line 1   Column 2917   Coefficient 69.29882813
   "010001010100110101", -- Line 1   Column 2918   Coefficient 69.30175781
   "010001010100111000", -- Line 1   Column 2919   Coefficient 69.30468750
   "010001010100111011", -- Line 1   Column 2920   Coefficient 69.30761719
   "010001010100111110", -- Line 1   Column 2921   Coefficient 69.31054688
   "010001010101000001", -- Line 1   Column 2922   Coefficient 69.31347656
   "010001010101000100", -- Line 1   Column 2923   Coefficient 69.31640625
   "010001010101000111", -- Line 1   Column 2924   Coefficient 69.31933594
   "010001010101001010", -- Line 1   Column 2925   Coefficient 69.32226563
   "010001010101001101", -- Line 1   Column 2926   Coefficient 69.32519531
   "010001010101010000", -- Line 1   Column 2927   Coefficient 69.32812500
   "010001010101010011", -- Line 1   Column 2928   Coefficient 69.33105469
   "010001010101010110", -- Line 1   Column 2929   Coefficient 69.33398438
   "010001010101011001", -- Line 1   Column 2930   Coefficient 69.33691406
   "010001010101011100", -- Line 1   Column 2931   Coefficient 69.33984375
   "010001010101100000", -- Line 1   Column 2932   Coefficient 69.34375000
   "010001010101100011", -- Line 1   Column 2933   Coefficient 69.34667969
   "010001010101100110", -- Line 1   Column 2934   Coefficient 69.34960938
   "010001010101101001", -- Line 1   Column 2935   Coefficient 69.35253906
   "010001010101101100", -- Line 1   Column 2936   Coefficient 69.35546875
   "010001010101101111", -- Line 1   Column 2937   Coefficient 69.35839844
   "010001010101110010", -- Line 1   Column 2938   Coefficient 69.36132813
   "010001010101110101", -- Line 1   Column 2939   Coefficient 69.36425781
   "010001010101111000", -- Line 1   Column 2940   Coefficient 69.36718750
   "010001010101111011", -- Line 1   Column 2941   Coefficient 69.37011719
   "010001010101111110", -- Line 1   Column 2942   Coefficient 69.37304688
   "010001010110000001", -- Line 1   Column 2943   Coefficient 69.37597656
   "010001010110000100", -- Line 1   Column 2944   Coefficient 69.37890625
   "010001010110000111", -- Line 1   Column 2945   Coefficient 69.38183594
   "010001010110001010", -- Line 1   Column 2946   Coefficient 69.38476563
   "010001010110001101", -- Line 1   Column 2947   Coefficient 69.38769531
   "010001010110010000", -- Line 1   Column 2948   Coefficient 69.39062500
   "010001010110010011", -- Line 1   Column 2949   Coefficient 69.39355469
   "010001010110010110", -- Line 1   Column 2950   Coefficient 69.39648438
   "010001010110011001", -- Line 1   Column 2951   Coefficient 69.39941406
   "010001010110011100", -- Line 1   Column 2952   Coefficient 69.40234375
   "010001010110011111", -- Line 1   Column 2953   Coefficient 69.40527344
   "010001010110100010", -- Line 1   Column 2954   Coefficient 69.40820313
   "010001010110100101", -- Line 1   Column 2955   Coefficient 69.41113281
   "010001010110101000", -- Line 1   Column 2956   Coefficient 69.41406250
   "010001010110101011", -- Line 1   Column 2957   Coefficient 69.41699219
   "010001010110101110", -- Line 1   Column 2958   Coefficient 69.41992188
   "010001010110110001", -- Line 1   Column 2959   Coefficient 69.42285156
   "010001010110110100", -- Line 1   Column 2960   Coefficient 69.42578125
   "010001010110110111", -- Line 1   Column 2961   Coefficient 69.42871094
   "010001010110111010", -- Line 1   Column 2962   Coefficient 69.43164063
   "010001010110111101", -- Line 1   Column 2963   Coefficient 69.43457031
   "010001010111000000", -- Line 1   Column 2964   Coefficient 69.43750000
   "010001010111000011", -- Line 1   Column 2965   Coefficient 69.44042969
   "010001010111000110", -- Line 1   Column 2966   Coefficient 69.44335938
   "010001010111001001", -- Line 1   Column 2967   Coefficient 69.44628906
   "010001010111001100", -- Line 1   Column 2968   Coefficient 69.44921875
   "010001010111001111", -- Line 1   Column 2969   Coefficient 69.45214844
   "010001010111010010", -- Line 1   Column 2970   Coefficient 69.45507813
   "010001010111010101", -- Line 1   Column 2971   Coefficient 69.45800781
   "010001010111011000", -- Line 1   Column 2972   Coefficient 69.46093750
   "010001010111011011", -- Line 1   Column 2973   Coefficient 69.46386719
   "010001010111011110", -- Line 1   Column 2974   Coefficient 69.46679688
   "010001010111100001", -- Line 1   Column 2975   Coefficient 69.46972656
   "010001010111100100", -- Line 1   Column 2976   Coefficient 69.47265625
   "010001010111100111", -- Line 1   Column 2977   Coefficient 69.47558594
   "010001010111101010", -- Line 1   Column 2978   Coefficient 69.47851563
   "010001010111101101", -- Line 1   Column 2979   Coefficient 69.48144531
   "010001010111110000", -- Line 1   Column 2980   Coefficient 69.48437500
   "010001010111110011", -- Line 1   Column 2981   Coefficient 69.48730469
   "010001010111110110", -- Line 1   Column 2982   Coefficient 69.49023438
   "010001010111111001", -- Line 1   Column 2983   Coefficient 69.49316406
   "010001010111111100", -- Line 1   Column 2984   Coefficient 69.49609375
   "010001010111111111", -- Line 1   Column 2985   Coefficient 69.49902344
   "010001011000000010", -- Line 1   Column 2986   Coefficient 69.50195313
   "010001011000000101", -- Line 1   Column 2987   Coefficient 69.50488281
   "010001011000001000", -- Line 1   Column 2988   Coefficient 69.50781250
   "010001011000001011", -- Line 1   Column 2989   Coefficient 69.51074219
   "010001011000001110", -- Line 1   Column 2990   Coefficient 69.51367188
   "010001011000010001", -- Line 1   Column 2991   Coefficient 69.51660156
   "010001011000010100", -- Line 1   Column 2992   Coefficient 69.51953125
   "010001011000010111", -- Line 1   Column 2993   Coefficient 69.52246094
   "010001011000011010", -- Line 1   Column 2994   Coefficient 69.52539063
   "010001011000011101", -- Line 1   Column 2995   Coefficient 69.52832031
   "010001011000100000", -- Line 1   Column 2996   Coefficient 69.53125000
   "010001011000100011", -- Line 1   Column 2997   Coefficient 69.53417969
   "010001011000100110", -- Line 1   Column 2998   Coefficient 69.53710938
   "010001011000101000", -- Line 1   Column 2999   Coefficient 69.53906250
   "010001011000101011", -- Line 1   Column 3000   Coefficient 69.54199219
   "010001011000101110", -- Line 1   Column 3001   Coefficient 69.54492188
   "010001011000110001", -- Line 1   Column 3002   Coefficient 69.54785156
   "010001011000110100", -- Line 1   Column 3003   Coefficient 69.55078125
   "010001011000110111", -- Line 1   Column 3004   Coefficient 69.55371094
   "010001011000111010", -- Line 1   Column 3005   Coefficient 69.55664063
   "010001011000111101", -- Line 1   Column 3006   Coefficient 69.55957031
   "010001011001000000", -- Line 1   Column 3007   Coefficient 69.56250000
   "010001011001000011", -- Line 1   Column 3008   Coefficient 69.56542969
   "010001011001000110", -- Line 1   Column 3009   Coefficient 69.56835938
   "010001011001001001", -- Line 1   Column 3010   Coefficient 69.57128906
   "010001011001001100", -- Line 1   Column 3011   Coefficient 69.57421875
   "010001011001001111", -- Line 1   Column 3012   Coefficient 69.57714844
   "010001011001010010", -- Line 1   Column 3013   Coefficient 69.58007813
   "010001011001010101", -- Line 1   Column 3014   Coefficient 69.58300781
   "010001011001011000", -- Line 1   Column 3015   Coefficient 69.58593750
   "010001011001011011", -- Line 1   Column 3016   Coefficient 69.58886719
   "010001011001011110", -- Line 1   Column 3017   Coefficient 69.59179688
   "010001011001100001", -- Line 1   Column 3018   Coefficient 69.59472656
   "010001011001100100", -- Line 1   Column 3019   Coefficient 69.59765625
   "010001011001100111", -- Line 1   Column 3020   Coefficient 69.60058594
   "010001011001101001", -- Line 1   Column 3021   Coefficient 69.60253906
   "010001011001101100", -- Line 1   Column 3022   Coefficient 69.60546875
   "010001011001101111", -- Line 1   Column 3023   Coefficient 69.60839844
   "010001011001110010", -- Line 1   Column 3024   Coefficient 69.61132813
   "010001011001110101", -- Line 1   Column 3025   Coefficient 69.61425781
   "010001011001111000", -- Line 1   Column 3026   Coefficient 69.61718750
   "010001011001111011", -- Line 1   Column 3027   Coefficient 69.62011719
   "010001011001111110", -- Line 1   Column 3028   Coefficient 69.62304688
   "010001011010000001", -- Line 1   Column 3029   Coefficient 69.62597656
   "010001011010000100", -- Line 1   Column 3030   Coefficient 69.62890625
   "010001011010000111", -- Line 1   Column 3031   Coefficient 69.63183594
   "010001011010001010", -- Line 1   Column 3032   Coefficient 69.63476563
   "010001011010001101", -- Line 1   Column 3033   Coefficient 69.63769531
   "010001011010010000", -- Line 1   Column 3034   Coefficient 69.64062500
   "010001011010010011", -- Line 1   Column 3035   Coefficient 69.64355469
   "010001011010010110", -- Line 1   Column 3036   Coefficient 69.64648438
   "010001011010011000", -- Line 1   Column 3037   Coefficient 69.64843750
   "010001011010011011", -- Line 1   Column 3038   Coefficient 69.65136719
   "010001011010011110", -- Line 1   Column 3039   Coefficient 69.65429688
   "010001011010100001", -- Line 1   Column 3040   Coefficient 69.65722656
   "010001011010100100", -- Line 1   Column 3041   Coefficient 69.66015625
   "010001011010100111", -- Line 1   Column 3042   Coefficient 69.66308594
   "010001011010101010", -- Line 1   Column 3043   Coefficient 69.66601563
   "010001011010101101", -- Line 1   Column 3044   Coefficient 69.66894531
   "010001011010110000", -- Line 1   Column 3045   Coefficient 69.67187500
   "010001011010110011", -- Line 1   Column 3046   Coefficient 69.67480469
   "010001011010110110", -- Line 1   Column 3047   Coefficient 69.67773438
   "010001011010111001", -- Line 1   Column 3048   Coefficient 69.68066406
   "010001011010111100", -- Line 1   Column 3049   Coefficient 69.68359375
   "010001011010111110", -- Line 1   Column 3050   Coefficient 69.68554688
   "010001011011000001", -- Line 1   Column 3051   Coefficient 69.68847656
   "010001011011000100", -- Line 1   Column 3052   Coefficient 69.69140625
   "010001011011000111", -- Line 1   Column 3053   Coefficient 69.69433594
   "010001011011001010", -- Line 1   Column 3054   Coefficient 69.69726563
   "010001011011001101", -- Line 1   Column 3055   Coefficient 69.70019531
   "010001011011010000", -- Line 1   Column 3056   Coefficient 69.70312500
   "010001011011010011", -- Line 1   Column 3057   Coefficient 69.70605469
   "010001011011010110", -- Line 1   Column 3058   Coefficient 69.70898438
   "010001011011011001", -- Line 1   Column 3059   Coefficient 69.71191406
   "010001011011011100", -- Line 1   Column 3060   Coefficient 69.71484375
   "010001011011011110", -- Line 1   Column 3061   Coefficient 69.71679688
   "010001011011100001", -- Line 1   Column 3062   Coefficient 69.71972656
   "010001011011100100", -- Line 1   Column 3063   Coefficient 69.72265625
   "010001011011100111", -- Line 1   Column 3064   Coefficient 69.72558594
   "010001011011101010", -- Line 1   Column 3065   Coefficient 69.72851563
   "010001011011101101", -- Line 1   Column 3066   Coefficient 69.73144531
   "010001011011110000", -- Line 1   Column 3067   Coefficient 69.73437500
   "010001011011110011", -- Line 1   Column 3068   Coefficient 69.73730469
   "010001011011110110", -- Line 1   Column 3069   Coefficient 69.74023438
   "010001011011111001", -- Line 1   Column 3070   Coefficient 69.74316406
   "010001011011111011", -- Line 1   Column 3071   Coefficient 69.74511719
   "010001011011111110", -- Line 1   Column 3072   Coefficient 69.74804688
   "010001011100000001", -- Line 1   Column 3073   Coefficient 69.75097656
   "010001011100000100", -- Line 1   Column 3074   Coefficient 69.75390625
   "010001011100000111", -- Line 1   Column 3075   Coefficient 69.75683594
   "010001011100001010", -- Line 1   Column 3076   Coefficient 69.75976563
   "010001011100001101", -- Line 1   Column 3077   Coefficient 69.76269531
   "010001011100010000", -- Line 1   Column 3078   Coefficient 69.76562500
   "010001011100010011", -- Line 1   Column 3079   Coefficient 69.76855469
   "010001011100010110", -- Line 1   Column 3080   Coefficient 69.77148438
   "010001011100011000", -- Line 1   Column 3081   Coefficient 69.77343750
   "010001011100011011", -- Line 1   Column 3082   Coefficient 69.77636719
   "010001011100011110", -- Line 1   Column 3083   Coefficient 69.77929688
   "010001011100100001", -- Line 1   Column 3084   Coefficient 69.78222656
   "010001011100100100", -- Line 1   Column 3085   Coefficient 69.78515625
   "010001011100100111", -- Line 1   Column 3086   Coefficient 69.78808594
   "010001011100101010", -- Line 1   Column 3087   Coefficient 69.79101563
   "010001011100101101", -- Line 1   Column 3088   Coefficient 69.79394531
   "010001011100101111", -- Line 1   Column 3089   Coefficient 69.79589844
   "010001011100110010", -- Line 1   Column 3090   Coefficient 69.79882813
   "010001011100110101", -- Line 1   Column 3091   Coefficient 69.80175781
   "010001011100111000", -- Line 1   Column 3092   Coefficient 69.80468750
   "010001011100111011", -- Line 1   Column 3093   Coefficient 69.80761719
   "010001011100111110", -- Line 1   Column 3094   Coefficient 69.81054688
   "010001011101000001", -- Line 1   Column 3095   Coefficient 69.81347656
   "010001011101000100", -- Line 1   Column 3096   Coefficient 69.81640625
   "010001011101000110", -- Line 1   Column 3097   Coefficient 69.81835938
   "010001011101001001", -- Line 1   Column 3098   Coefficient 69.82128906
   "010001011101001100", -- Line 1   Column 3099   Coefficient 69.82421875
   "010001011101001111", -- Line 1   Column 3100   Coefficient 69.82714844
   "010001011101010010", -- Line 1   Column 3101   Coefficient 69.83007813
   "010001011101010101", -- Line 1   Column 3102   Coefficient 69.83300781
   "010001011101011000", -- Line 1   Column 3103   Coefficient 69.83593750
   "010001011101011011", -- Line 1   Column 3104   Coefficient 69.83886719
   "010001011101011101", -- Line 1   Column 3105   Coefficient 69.84082031
   "010001011101100000", -- Line 1   Column 3106   Coefficient 69.84375000
   "010001011101100011", -- Line 1   Column 3107   Coefficient 69.84667969
   "010001011101100110", -- Line 1   Column 3108   Coefficient 69.84960938
   "010001011101101001", -- Line 1   Column 3109   Coefficient 69.85253906
   "010001011101101100", -- Line 1   Column 3110   Coefficient 69.85546875
   "010001011101101111", -- Line 1   Column 3111   Coefficient 69.85839844
   "010001011101110001", -- Line 1   Column 3112   Coefficient 69.86035156
   "010001011101110100", -- Line 1   Column 3113   Coefficient 69.86328125
   "010001011101110111", -- Line 1   Column 3114   Coefficient 69.86621094
   "010001011101111010", -- Line 1   Column 3115   Coefficient 69.86914063
   "010001011101111101", -- Line 1   Column 3116   Coefficient 69.87207031
   "010001011110000000", -- Line 1   Column 3117   Coefficient 69.87500000
   "010001011110000011", -- Line 1   Column 3118   Coefficient 69.87792969
   "010001011110000101", -- Line 1   Column 3119   Coefficient 69.87988281
   "010001011110001000", -- Line 1   Column 3120   Coefficient 69.88281250
   "010001011110001011", -- Line 1   Column 3121   Coefficient 69.88574219
   "010001011110001110", -- Line 1   Column 3122   Coefficient 69.88867188
   "010001011110010001", -- Line 1   Column 3123   Coefficient 69.89160156
   "010001011110010100", -- Line 1   Column 3124   Coefficient 69.89453125
   "010001011110010111", -- Line 1   Column 3125   Coefficient 69.89746094
   "010001011110011001", -- Line 1   Column 3126   Coefficient 69.89941406
   "010001011110011100", -- Line 1   Column 3127   Coefficient 69.90234375
   "010001011110011111", -- Line 1   Column 3128   Coefficient 69.90527344
   "010001011110100010", -- Line 1   Column 3129   Coefficient 69.90820313
   "010001011110100101", -- Line 1   Column 3130   Coefficient 69.91113281
   "010001011110101000", -- Line 1   Column 3131   Coefficient 69.91406250
   "010001011110101010", -- Line 1   Column 3132   Coefficient 69.91601563
   "010001011110101101", -- Line 1   Column 3133   Coefficient 69.91894531
   "010001011110110000", -- Line 1   Column 3134   Coefficient 69.92187500
   "010001011110110011", -- Line 1   Column 3135   Coefficient 69.92480469
   "010001011110110110", -- Line 1   Column 3136   Coefficient 69.92773438
   "010001011110111001", -- Line 1   Column 3137   Coefficient 69.93066406
   "010001011110111011", -- Line 1   Column 3138   Coefficient 69.93261719
   "010001011110111110", -- Line 1   Column 3139   Coefficient 69.93554688
   "010001011111000001", -- Line 1   Column 3140   Coefficient 69.93847656
   "010001011111000100", -- Line 1   Column 3141   Coefficient 69.94140625
   "010001011111000111", -- Line 1   Column 3142   Coefficient 69.94433594
   "010001011111001010", -- Line 1   Column 3143   Coefficient 69.94726563
   "010001011111001100", -- Line 1   Column 3144   Coefficient 69.94921875
   "010001011111001111", -- Line 1   Column 3145   Coefficient 69.95214844
   "010001011111010010", -- Line 1   Column 3146   Coefficient 69.95507813
   "010001011111010101", -- Line 1   Column 3147   Coefficient 69.95800781
   "010001011111011000", -- Line 1   Column 3148   Coefficient 69.96093750
   "010001011111011011", -- Line 1   Column 3149   Coefficient 69.96386719
   "010001011111011101", -- Line 1   Column 3150   Coefficient 69.96582031
   "010001011111100000", -- Line 1   Column 3151   Coefficient 69.96875000
   "010001011111100011", -- Line 1   Column 3152   Coefficient 69.97167969
   "010001011111100110", -- Line 1   Column 3153   Coefficient 69.97460938
   "010001011111101001", -- Line 1   Column 3154   Coefficient 69.97753906
   "010001011111101100", -- Line 1   Column 3155   Coefficient 69.98046875
   "010001011111101110", -- Line 1   Column 3156   Coefficient 69.98242188
   "010001011111110001", -- Line 1   Column 3157   Coefficient 69.98535156
   "010001011111110100", -- Line 1   Column 3158   Coefficient 69.98828125
   "010001011111110111", -- Line 1   Column 3159   Coefficient 69.99121094
   "010001011111111010", -- Line 1   Column 3160   Coefficient 69.99414063
   "010001011111111100", -- Line 1   Column 3161   Coefficient 69.99609375
   "010001011111111111", -- Line 1   Column 3162   Coefficient 69.99902344
   "010001100000000010", -- Line 1   Column 3163   Coefficient 70.00195313
   "010001100000000101", -- Line 1   Column 3164   Coefficient 70.00488281
   "010001100000001000", -- Line 1   Column 3165   Coefficient 70.00781250
   "010001100000001010", -- Line 1   Column 3166   Coefficient 70.00976563
   "010001100000001101", -- Line 1   Column 3167   Coefficient 70.01269531
   "010001100000010000", -- Line 1   Column 3168   Coefficient 70.01562500
   "010001100000010011", -- Line 1   Column 3169   Coefficient 70.01855469
   "010001100000010110", -- Line 1   Column 3170   Coefficient 70.02148438
   "010001100000011000", -- Line 1   Column 3171   Coefficient 70.02343750
   "010001100000011011", -- Line 1   Column 3172   Coefficient 70.02636719
   "010001100000011110", -- Line 1   Column 3173   Coefficient 70.02929688
   "010001100000100001", -- Line 1   Column 3174   Coefficient 70.03222656
   "010001100000100100", -- Line 1   Column 3175   Coefficient 70.03515625
   "010001100000100111", -- Line 1   Column 3176   Coefficient 70.03808594
   "010001100000101001", -- Line 1   Column 3177   Coefficient 70.04003906
   "010001100000101100", -- Line 1   Column 3178   Coefficient 70.04296875
   "010001100000101111", -- Line 1   Column 3179   Coefficient 70.04589844
   "010001100000110010", -- Line 1   Column 3180   Coefficient 70.04882813
   "010001100000110101", -- Line 1   Column 3181   Coefficient 70.05175781
   "010001100000110111", -- Line 1   Column 3182   Coefficient 70.05371094
   "010001100000111010", -- Line 1   Column 3183   Coefficient 70.05664063
   "010001100000111101", -- Line 1   Column 3184   Coefficient 70.05957031
   "010001100001000000", -- Line 1   Column 3185   Coefficient 70.06250000
   "010001100001000010", -- Line 1   Column 3186   Coefficient 70.06445313
   "010001100001000101", -- Line 1   Column 3187   Coefficient 70.06738281
   "010001100001001000", -- Line 1   Column 3188   Coefficient 70.07031250
   "010001100001001011", -- Line 1   Column 3189   Coefficient 70.07324219
   "010001100001001110", -- Line 1   Column 3190   Coefficient 70.07617188
   "010001100001010000", -- Line 1   Column 3191   Coefficient 70.07812500
   "010001100001010011", -- Line 1   Column 3192   Coefficient 70.08105469
   "010001100001010110", -- Line 1   Column 3193   Coefficient 70.08398438
   "010001100001011001", -- Line 1   Column 3194   Coefficient 70.08691406
   "010001100001011100", -- Line 1   Column 3195   Coefficient 70.08984375
   "010001100001011110", -- Line 1   Column 3196   Coefficient 70.09179688
   "010001100001100001", -- Line 1   Column 3197   Coefficient 70.09472656
   "010001100001100100", -- Line 1   Column 3198   Coefficient 70.09765625
   "010001100001100111", -- Line 1   Column 3199   Coefficient 70.10058594
   "010001100001101001", -- Line 1   Column 3200   Coefficient 70.10253906
   "010001100001101100", -- Line 1   Column 3201   Coefficient 70.10546875
   "010001100001101111", -- Line 1   Column 3202   Coefficient 70.10839844
   "010001100001110010", -- Line 1   Column 3203   Coefficient 70.11132813
   "010001100001110101", -- Line 1   Column 3204   Coefficient 70.11425781
   "010001100001110111", -- Line 1   Column 3205   Coefficient 70.11621094
   "010001100001111010", -- Line 1   Column 3206   Coefficient 70.11914063
   "010001100001111101", -- Line 1   Column 3207   Coefficient 70.12207031
   "010001100010000000", -- Line 1   Column 3208   Coefficient 70.12500000
   "010001100010000010", -- Line 1   Column 3209   Coefficient 70.12695313
   "010001100010000101", -- Line 1   Column 3210   Coefficient 70.12988281
   "010001100010001000", -- Line 1   Column 3211   Coefficient 70.13281250
   "010001100010001011", -- Line 1   Column 3212   Coefficient 70.13574219
   "010001100010001110", -- Line 1   Column 3213   Coefficient 70.13867188
   "010001100010010000", -- Line 1   Column 3214   Coefficient 70.14062500
   "010001100010010011", -- Line 1   Column 3215   Coefficient 70.14355469
   "010001100010010110", -- Line 1   Column 3216   Coefficient 70.14648438
   "010001100010011001", -- Line 1   Column 3217   Coefficient 70.14941406
   "010001100010011011", -- Line 1   Column 3218   Coefficient 70.15136719
   "010001100010011110", -- Line 1   Column 3219   Coefficient 70.15429688
   "010001100010100001", -- Line 1   Column 3220   Coefficient 70.15722656
   "010001100010100100", -- Line 1   Column 3221   Coefficient 70.16015625
   "010001100010100110", -- Line 1   Column 3222   Coefficient 70.16210938
   "010001100010101001", -- Line 1   Column 3223   Coefficient 70.16503906
   "010001100010101100", -- Line 1   Column 3224   Coefficient 70.16796875
   "010001100010101111", -- Line 1   Column 3225   Coefficient 70.17089844
   "010001100010110001", -- Line 1   Column 3226   Coefficient 70.17285156
   "010001100010110100", -- Line 1   Column 3227   Coefficient 70.17578125
   "010001100010110111", -- Line 1   Column 3228   Coefficient 70.17871094
   "010001100010111010", -- Line 1   Column 3229   Coefficient 70.18164063
   "010001100010111100", -- Line 1   Column 3230   Coefficient 70.18359375
   "010001100010111111", -- Line 1   Column 3231   Coefficient 70.18652344
   "010001100011000010", -- Line 1   Column 3232   Coefficient 70.18945313
   "010001100011000101", -- Line 1   Column 3233   Coefficient 70.19238281
   "010001100011000111", -- Line 1   Column 3234   Coefficient 70.19433594
   "010001100011001010", -- Line 1   Column 3235   Coefficient 70.19726563
   "010001100011001101", -- Line 1   Column 3236   Coefficient 70.20019531
   "010001100011010000", -- Line 1   Column 3237   Coefficient 70.20312500
   "010001100011010010", -- Line 1   Column 3238   Coefficient 70.20507813
   "010001100011010101", -- Line 1   Column 3239   Coefficient 70.20800781
   "010001100011011000", -- Line 1   Column 3240   Coefficient 70.21093750
   "010001100011011011", -- Line 1   Column 3241   Coefficient 70.21386719
   "010001100011011101", -- Line 1   Column 3242   Coefficient 70.21582031
   "010001100011100000", -- Line 1   Column 3243   Coefficient 70.21875000
   "010001100011100011", -- Line 1   Column 3244   Coefficient 70.22167969
   "010001100011100110", -- Line 1   Column 3245   Coefficient 70.22460938
   "010001100011101000", -- Line 1   Column 3246   Coefficient 70.22656250
   "010001100011101011", -- Line 1   Column 3247   Coefficient 70.22949219
   "010001100011101110", -- Line 1   Column 3248   Coefficient 70.23242188
   "010001100011110001", -- Line 1   Column 3249   Coefficient 70.23535156
   "010001100011110011", -- Line 1   Column 3250   Coefficient 70.23730469
   "010001100011110110", -- Line 1   Column 3251   Coefficient 70.24023438
   "010001100011111001", -- Line 1   Column 3252   Coefficient 70.24316406
   "010001100011111100", -- Line 1   Column 3253   Coefficient 70.24609375
   "010001100011111110", -- Line 1   Column 3254   Coefficient 70.24804688
   "010001100100000001", -- Line 1   Column 3255   Coefficient 70.25097656
   "010001100100000100", -- Line 1   Column 3256   Coefficient 70.25390625
   "010001100100000111", -- Line 1   Column 3257   Coefficient 70.25683594
   "010001100100001001", -- Line 1   Column 3258   Coefficient 70.25878906
   "010001100100001100", -- Line 1   Column 3259   Coefficient 70.26171875
   "010001100100001111", -- Line 1   Column 3260   Coefficient 70.26464844
   "010001100100010001", -- Line 1   Column 3261   Coefficient 70.26660156
   "010001100100010100", -- Line 1   Column 3262   Coefficient 70.26953125
   "010001100100010111", -- Line 1   Column 3263   Coefficient 70.27246094
   "010001100100011010", -- Line 1   Column 3264   Coefficient 70.27539063
   "010001100100011100", -- Line 1   Column 3265   Coefficient 70.27734375
   "010001100100011111", -- Line 1   Column 3266   Coefficient 70.28027344
   "010001100100100010", -- Line 1   Column 3267   Coefficient 70.28320313
   "010001100100100100", -- Line 1   Column 3268   Coefficient 70.28515625
   "010001100100100111", -- Line 1   Column 3269   Coefficient 70.28808594
   "010001100100101010", -- Line 1   Column 3270   Coefficient 70.29101563
   "010001100100101101", -- Line 1   Column 3271   Coefficient 70.29394531
   "010001100100101111", -- Line 1   Column 3272   Coefficient 70.29589844
   "010001100100110010", -- Line 1   Column 3273   Coefficient 70.29882813
   "010001100100110101", -- Line 1   Column 3274   Coefficient 70.30175781
   "010001100100111000", -- Line 1   Column 3275   Coefficient 70.30468750
   "010001100100111010", -- Line 1   Column 3276   Coefficient 70.30664063
   "010001100100111101", -- Line 1   Column 3277   Coefficient 70.30957031
   "010001100101000000", -- Line 1   Column 3278   Coefficient 70.31250000
   "010001100101000010", -- Line 1   Column 3279   Coefficient 70.31445313
   "010001100101000101", -- Line 1   Column 3280   Coefficient 70.31738281
   "010001100101001000", -- Line 1   Column 3281   Coefficient 70.32031250
   "010001100101001011", -- Line 1   Column 3282   Coefficient 70.32324219
   "010001100101001101", -- Line 1   Column 3283   Coefficient 70.32519531
   "010001100101010000", -- Line 1   Column 3284   Coefficient 70.32812500
   "010001100101010011", -- Line 1   Column 3285   Coefficient 70.33105469
   "010001100101010101", -- Line 1   Column 3286   Coefficient 70.33300781
   "010001100101011000", -- Line 1   Column 3287   Coefficient 70.33593750
   "010001100101011011", -- Line 1   Column 3288   Coefficient 70.33886719
   "010001100101011101", -- Line 1   Column 3289   Coefficient 70.34082031
   "010001100101100000", -- Line 1   Column 3290   Coefficient 70.34375000
   "010001100101100011", -- Line 1   Column 3291   Coefficient 70.34667969
   "010001100101100110", -- Line 1   Column 3292   Coefficient 70.34960938
   "010001100101101000", -- Line 1   Column 3293   Coefficient 70.35156250
   "010001100101101011", -- Line 1   Column 3294   Coefficient 70.35449219
   "010001100101101110", -- Line 1   Column 3295   Coefficient 70.35742188
   "010001100101110000", -- Line 1   Column 3296   Coefficient 70.35937500
   "010001100101110011", -- Line 1   Column 3297   Coefficient 70.36230469
   "010001100101110110", -- Line 1   Column 3298   Coefficient 70.36523438
   "010001100101111000", -- Line 1   Column 3299   Coefficient 70.36718750
   "010001100101111011", -- Line 1   Column 3300   Coefficient 70.37011719
   "010001100101111110", -- Line 1   Column 3301   Coefficient 70.37304688
   "010001100110000001", -- Line 1   Column 3302   Coefficient 70.37597656
   "010001100110000011", -- Line 1   Column 3303   Coefficient 70.37792969
   "010001100110000110", -- Line 1   Column 3304   Coefficient 70.38085938
   "010001100110001001", -- Line 1   Column 3305   Coefficient 70.38378906
   "010001100110001011", -- Line 1   Column 3306   Coefficient 70.38574219
   "010001100110001110", -- Line 1   Column 3307   Coefficient 70.38867188
   "010001100110010001", -- Line 1   Column 3308   Coefficient 70.39160156
   "010001100110010011", -- Line 1   Column 3309   Coefficient 70.39355469
   "010001100110010110", -- Line 1   Column 3310   Coefficient 70.39648438
   "010001100110011001", -- Line 1   Column 3311   Coefficient 70.39941406
   "010001100110011011", -- Line 1   Column 3312   Coefficient 70.40136719
   "010001100110011110", -- Line 1   Column 3313   Coefficient 70.40429688
   "010001100110100001", -- Line 1   Column 3314   Coefficient 70.40722656
   "010001100110100100", -- Line 1   Column 3315   Coefficient 70.41015625
   "010001100110100110", -- Line 1   Column 3316   Coefficient 70.41210938
   "010001100110101001", -- Line 1   Column 3317   Coefficient 70.41503906
   "010001100110101100", -- Line 1   Column 3318   Coefficient 70.41796875
   "010001100110101110", -- Line 1   Column 3319   Coefficient 70.41992188
   "010001100110110001", -- Line 1   Column 3320   Coefficient 70.42285156
   "010001100110110100", -- Line 1   Column 3321   Coefficient 70.42578125
   "010001100110110110", -- Line 1   Column 3322   Coefficient 70.42773438
   "010001100110111001", -- Line 1   Column 3323   Coefficient 70.43066406
   "010001100110111100", -- Line 1   Column 3324   Coefficient 70.43359375
   "010001100110111110", -- Line 1   Column 3325   Coefficient 70.43554688
   "010001100111000001", -- Line 1   Column 3326   Coefficient 70.43847656
   "010001100111000100", -- Line 1   Column 3327   Coefficient 70.44140625
   "010001100111000110", -- Line 1   Column 3328   Coefficient 70.44335938
   "010001100111001001", -- Line 1   Column 3329   Coefficient 70.44628906
   "010001100111001100", -- Line 1   Column 3330   Coefficient 70.44921875
   "010001100111001110", -- Line 1   Column 3331   Coefficient 70.45117188
   "010001100111010001", -- Line 1   Column 3332   Coefficient 70.45410156
   "010001100111010100", -- Line 1   Column 3333   Coefficient 70.45703125
   "010001100111010110", -- Line 1   Column 3334   Coefficient 70.45898438
   "010001100111011001", -- Line 1   Column 3335   Coefficient 70.46191406
   "010001100111011100", -- Line 1   Column 3336   Coefficient 70.46484375
   "010001100111011110", -- Line 1   Column 3337   Coefficient 70.46679688
   "010001100111100001", -- Line 1   Column 3338   Coefficient 70.46972656
   "010001100111100100", -- Line 1   Column 3339   Coefficient 70.47265625
   "010001100111100110", -- Line 1   Column 3340   Coefficient 70.47460938
   "010001100111101001", -- Line 1   Column 3341   Coefficient 70.47753906
   "010001100111101100", -- Line 1   Column 3342   Coefficient 70.48046875
   "010001100111101110", -- Line 1   Column 3343   Coefficient 70.48242188
   "010001100111110001", -- Line 1   Column 3344   Coefficient 70.48535156
   "010001100111110100", -- Line 1   Column 3345   Coefficient 70.48828125
   "010001100111110110", -- Line 1   Column 3346   Coefficient 70.49023438
   "010001100111111001", -- Line 1   Column 3347   Coefficient 70.49316406
   "010001100111111100", -- Line 1   Column 3348   Coefficient 70.49609375
   "010001100111111110", -- Line 1   Column 3349   Coefficient 70.49804688
   "010001101000000001", -- Line 1   Column 3350   Coefficient 70.50097656
   "010001101000000100", -- Line 1   Column 3351   Coefficient 70.50390625
   "010001101000000110", -- Line 1   Column 3352   Coefficient 70.50585938
   "010001101000001001", -- Line 1   Column 3353   Coefficient 70.50878906
   "010001101000001100", -- Line 1   Column 3354   Coefficient 70.51171875
   "010001101000001110", -- Line 1   Column 3355   Coefficient 70.51367188
   "010001101000010001", -- Line 1   Column 3356   Coefficient 70.51660156
   "010001101000010011", -- Line 1   Column 3357   Coefficient 70.51855469
   "010001101000010110", -- Line 1   Column 3358   Coefficient 70.52148438
   "010001101000011001", -- Line 1   Column 3359   Coefficient 70.52441406
   "010001101000011011", -- Line 1   Column 3360   Coefficient 70.52636719
   "010001101000011110", -- Line 1   Column 3361   Coefficient 70.52929688
   "010001101000100001", -- Line 1   Column 3362   Coefficient 70.53222656
   "010001101000100011", -- Line 1   Column 3363   Coefficient 70.53417969
   "010001101000100110", -- Line 1   Column 3364   Coefficient 70.53710938
   "010001101000101001", -- Line 1   Column 3365   Coefficient 70.54003906
   "010001101000101011", -- Line 1   Column 3366   Coefficient 70.54199219
   "010001101000101110", -- Line 1   Column 3367   Coefficient 70.54492188
   "010001101000110001", -- Line 1   Column 3368   Coefficient 70.54785156
   "010001101000110011", -- Line 1   Column 3369   Coefficient 70.54980469
   "010001101000110110", -- Line 1   Column 3370   Coefficient 70.55273438
   "010001101000111000", -- Line 1   Column 3371   Coefficient 70.55468750
   "010001101000111011", -- Line 1   Column 3372   Coefficient 70.55761719
   "010001101000111110", -- Line 1   Column 3373   Coefficient 70.56054688
   "010001101001000000", -- Line 1   Column 3374   Coefficient 70.56250000
   "010001101001000011", -- Line 1   Column 3375   Coefficient 70.56542969
   "010001101001000110", -- Line 1   Column 3376   Coefficient 70.56835938
   "010001101001001000", -- Line 1   Column 3377   Coefficient 70.57031250
   "010001101001001011", -- Line 1   Column 3378   Coefficient 70.57324219
   "010001101001001110", -- Line 1   Column 3379   Coefficient 70.57617188
   "010001101001010000", -- Line 1   Column 3380   Coefficient 70.57812500
   "010001101001010011", -- Line 1   Column 3381   Coefficient 70.58105469
   "010001101001010101", -- Line 1   Column 3382   Coefficient 70.58300781
   "010001101001011000", -- Line 1   Column 3383   Coefficient 70.58593750
   "010001101001011011", -- Line 1   Column 3384   Coefficient 70.58886719
   "010001101001011101", -- Line 1   Column 3385   Coefficient 70.59082031
   "010001101001100000", -- Line 1   Column 3386   Coefficient 70.59375000
   "010001101001100011", -- Line 1   Column 3387   Coefficient 70.59667969
   "010001101001100101", -- Line 1   Column 3388   Coefficient 70.59863281
   "010001101001101000", -- Line 1   Column 3389   Coefficient 70.60156250
   "010001101001101010", -- Line 1   Column 3390   Coefficient 70.60351563
   "010001101001101101", -- Line 1   Column 3391   Coefficient 70.60644531
   "010001101001110000", -- Line 1   Column 3392   Coefficient 70.60937500
   "010001101001110010", -- Line 1   Column 3393   Coefficient 70.61132813
   "010001101001110101", -- Line 1   Column 3394   Coefficient 70.61425781
   "010001101001111000", -- Line 1   Column 3395   Coefficient 70.61718750
   "010001101001111010", -- Line 1   Column 3396   Coefficient 70.61914063
   "010001101001111101", -- Line 1   Column 3397   Coefficient 70.62207031
   "010001101001111111", -- Line 1   Column 3398   Coefficient 70.62402344
   "010001101010000010", -- Line 1   Column 3399   Coefficient 70.62695313
   "010001101010000101", -- Line 1   Column 3400   Coefficient 70.62988281
   "010001101010000111", -- Line 1   Column 3401   Coefficient 70.63183594
   "010001101010001010", -- Line 1   Column 3402   Coefficient 70.63476563
   "010001101010001101", -- Line 1   Column 3403   Coefficient 70.63769531
   "010001101010001111", -- Line 1   Column 3404   Coefficient 70.63964844
   "010001101010010010", -- Line 1   Column 3405   Coefficient 70.64257813
   "010001101010010100", -- Line 1   Column 3406   Coefficient 70.64453125
   "010001101010010111", -- Line 1   Column 3407   Coefficient 70.64746094
   "010001101010011010", -- Line 1   Column 3408   Coefficient 70.65039063
   "010001101010011100", -- Line 1   Column 3409   Coefficient 70.65234375
   "010001101010011111", -- Line 1   Column 3410   Coefficient 70.65527344
   "010001101010100001", -- Line 1   Column 3411   Coefficient 70.65722656
   "010001101010100100", -- Line 1   Column 3412   Coefficient 70.66015625
   "010001101010100111", -- Line 1   Column 3413   Coefficient 70.66308594
   "010001101010101001", -- Line 1   Column 3414   Coefficient 70.66503906
   "010001101010101100", -- Line 1   Column 3415   Coefficient 70.66796875
   "010001101010101110", -- Line 1   Column 3416   Coefficient 70.66992188
   "010001101010110001", -- Line 1   Column 3417   Coefficient 70.67285156
   "010001101010110100", -- Line 1   Column 3418   Coefficient 70.67578125
   "010001101010110110", -- Line 1   Column 3419   Coefficient 70.67773438
   "010001101010111001", -- Line 1   Column 3420   Coefficient 70.68066406
   "010001101010111011", -- Line 1   Column 3421   Coefficient 70.68261719
   "010001101010111110", -- Line 1   Column 3422   Coefficient 70.68554688
   "010001101011000001", -- Line 1   Column 3423   Coefficient 70.68847656
   "010001101011000011", -- Line 1   Column 3424   Coefficient 70.69042969
   "010001101011000110", -- Line 1   Column 3425   Coefficient 70.69335938
   "010001101011001000", -- Line 1   Column 3426   Coefficient 70.69531250
   "010001101011001011", -- Line 1   Column 3427   Coefficient 70.69824219
   "010001101011001110", -- Line 1   Column 3428   Coefficient 70.70117188
   "010001101011010000", -- Line 1   Column 3429   Coefficient 70.70312500
   "010001101011010011", -- Line 1   Column 3430   Coefficient 70.70605469
   "010001101011010101", -- Line 1   Column 3431   Coefficient 70.70800781
   "010001101011011000", -- Line 1   Column 3432   Coefficient 70.71093750
   "010001101011011011", -- Line 1   Column 3433   Coefficient 70.71386719
   "010001101011011101", -- Line 1   Column 3434   Coefficient 70.71582031
   "010001101011100000", -- Line 1   Column 3435   Coefficient 70.71875000
   "010001101011100010", -- Line 1   Column 3436   Coefficient 70.72070313
   "010001101011100101", -- Line 1   Column 3437   Coefficient 70.72363281
   "010001101011101000", -- Line 1   Column 3438   Coefficient 70.72656250
   "010001101011101010", -- Line 1   Column 3439   Coefficient 70.72851563
   "010001101011101101", -- Line 1   Column 3440   Coefficient 70.73144531
   "010001101011101111", -- Line 1   Column 3441   Coefficient 70.73339844
   "010001101011110010", -- Line 1   Column 3442   Coefficient 70.73632813
   "010001101011110100", -- Line 1   Column 3443   Coefficient 70.73828125
   "010001101011110111", -- Line 1   Column 3444   Coefficient 70.74121094
   "010001101011111010", -- Line 1   Column 3445   Coefficient 70.74414063
   "010001101011111100", -- Line 1   Column 3446   Coefficient 70.74609375
   "010001101011111111", -- Line 1   Column 3447   Coefficient 70.74902344
   "010001101100000001", -- Line 1   Column 3448   Coefficient 70.75097656
   "010001101100000100", -- Line 1   Column 3449   Coefficient 70.75390625
   "010001101100000111", -- Line 1   Column 3450   Coefficient 70.75683594
   "010001101100001001", -- Line 1   Column 3451   Coefficient 70.75878906
   "010001101100001100", -- Line 1   Column 3452   Coefficient 70.76171875
   "010001101100001110", -- Line 1   Column 3453   Coefficient 70.76367188
   "010001101100010001", -- Line 1   Column 3454   Coefficient 70.76660156
   "010001101100010011", -- Line 1   Column 3455   Coefficient 70.76855469
   "010001101100010110", -- Line 1   Column 3456   Coefficient 70.77148438
   "010001101100011001", -- Line 1   Column 3457   Coefficient 70.77441406
   "010001101100011011", -- Line 1   Column 3458   Coefficient 70.77636719
   "010001101100011110", -- Line 1   Column 3459   Coefficient 70.77929688
   "010001101100100000", -- Line 1   Column 3460   Coefficient 70.78125000
   "010001101100100011", -- Line 1   Column 3461   Coefficient 70.78417969
   "010001101100100101", -- Line 1   Column 3462   Coefficient 70.78613281
   "010001101100101000", -- Line 1   Column 3463   Coefficient 70.78906250
   "010001101100101011", -- Line 1   Column 3464   Coefficient 70.79199219
   "010001101100101101", -- Line 1   Column 3465   Coefficient 70.79394531
   "010001101100110000", -- Line 1   Column 3466   Coefficient 70.79687500
   "010001101100110010", -- Line 1   Column 3467   Coefficient 70.79882813
   "010001101100110101", -- Line 1   Column 3468   Coefficient 70.80175781
   "010001101100110111", -- Line 1   Column 3469   Coefficient 70.80371094
   "010001101100111010", -- Line 1   Column 3470   Coefficient 70.80664063
   "010001101100111101", -- Line 1   Column 3471   Coefficient 70.80957031
   "010001101100111111", -- Line 1   Column 3472   Coefficient 70.81152344
   "010001101101000010", -- Line 1   Column 3473   Coefficient 70.81445313
   "010001101101000100", -- Line 1   Column 3474   Coefficient 70.81640625
   "010001101101000111", -- Line 1   Column 3475   Coefficient 70.81933594
   "010001101101001001", -- Line 1   Column 3476   Coefficient 70.82128906
   "010001101101001100", -- Line 1   Column 3477   Coefficient 70.82421875
   "010001101101001110", -- Line 1   Column 3478   Coefficient 70.82617188
   "010001101101010001", -- Line 1   Column 3479   Coefficient 70.82910156
   "010001101101010100", -- Line 1   Column 3480   Coefficient 70.83203125
   "010001101101010110", -- Line 1   Column 3481   Coefficient 70.83398438
   "010001101101011001", -- Line 1   Column 3482   Coefficient 70.83691406
   "010001101101011011", -- Line 1   Column 3483   Coefficient 70.83886719
   "010001101101011110", -- Line 1   Column 3484   Coefficient 70.84179688
   "010001101101100000", -- Line 1   Column 3485   Coefficient 70.84375000
   "010001101101100011", -- Line 1   Column 3486   Coefficient 70.84667969
   "010001101101100101", -- Line 1   Column 3487   Coefficient 70.84863281
   "010001101101101000", -- Line 1   Column 3488   Coefficient 70.85156250
   "010001101101101011", -- Line 1   Column 3489   Coefficient 70.85449219
   "010001101101101101", -- Line 1   Column 3490   Coefficient 70.85644531
   "010001101101110000", -- Line 1   Column 3491   Coefficient 70.85937500
   "010001101101110010", -- Line 1   Column 3492   Coefficient 70.86132813
   "010001101101110101", -- Line 1   Column 3493   Coefficient 70.86425781
   "010001101101110111", -- Line 1   Column 3494   Coefficient 70.86621094
   "010001101101111010", -- Line 1   Column 3495   Coefficient 70.86914063
   "010001101101111100", -- Line 1   Column 3496   Coefficient 70.87109375
   "010001101101111111", -- Line 1   Column 3497   Coefficient 70.87402344
   "010001101110000001", -- Line 1   Column 3498   Coefficient 70.87597656
   "010001101110000100", -- Line 1   Column 3499   Coefficient 70.87890625
   "010001101110000111", -- Line 1   Column 3500   Coefficient 70.88183594
   "010001101110001001", -- Line 1   Column 3501   Coefficient 70.88378906
   "010001101110001100", -- Line 1   Column 3502   Coefficient 70.88671875
   "010001101110001110", -- Line 1   Column 3503   Coefficient 70.88867188
   "010001101110010001", -- Line 1   Column 3504   Coefficient 70.89160156
   "010001101110010011", -- Line 1   Column 3505   Coefficient 70.89355469
   "010001101110010110", -- Line 1   Column 3506   Coefficient 70.89648438
   "010001101110011000", -- Line 1   Column 3507   Coefficient 70.89843750
   "010001101110011011", -- Line 1   Column 3508   Coefficient 70.90136719
   "010001101110011101", -- Line 1   Column 3509   Coefficient 70.90332031
   "010001101110100000", -- Line 1   Column 3510   Coefficient 70.90625000
   "010001101110100010", -- Line 1   Column 3511   Coefficient 70.90820313
   "010001101110100101", -- Line 1   Column 3512   Coefficient 70.91113281
   "010001101110100111", -- Line 1   Column 3513   Coefficient 70.91308594
   "010001101110101010", -- Line 1   Column 3514   Coefficient 70.91601563
   "010001101110101101", -- Line 1   Column 3515   Coefficient 70.91894531
   "010001101110101111", -- Line 1   Column 3516   Coefficient 70.92089844
   "010001101110110010", -- Line 1   Column 3517   Coefficient 70.92382813
   "010001101110110100", -- Line 1   Column 3518   Coefficient 70.92578125
   "010001101110110111", -- Line 1   Column 3519   Coefficient 70.92871094
   "010001101110111001", -- Line 1   Column 3520   Coefficient 70.93066406
   "010001101110111100", -- Line 1   Column 3521   Coefficient 70.93359375
   "010001101110111110", -- Line 1   Column 3522   Coefficient 70.93554688
   "010001101111000001", -- Line 1   Column 3523   Coefficient 70.93847656
   "010001101111000011", -- Line 1   Column 3524   Coefficient 70.94042969
   "010001101111000110", -- Line 1   Column 3525   Coefficient 70.94335938
   "010001101111001000", -- Line 1   Column 3526   Coefficient 70.94531250
   "010001101111001011", -- Line 1   Column 3527   Coefficient 70.94824219
   "010001101111001101", -- Line 1   Column 3528   Coefficient 70.95019531
   "010001101111010000", -- Line 1   Column 3529   Coefficient 70.95312500
   "010001101111010010", -- Line 1   Column 3530   Coefficient 70.95507813
   "010001101111010101", -- Line 1   Column 3531   Coefficient 70.95800781
   "010001101111010111", -- Line 1   Column 3532   Coefficient 70.95996094
   "010001101111011010", -- Line 1   Column 3533   Coefficient 70.96289063
   "010001101111011100", -- Line 1   Column 3534   Coefficient 70.96484375
   "010001101111011111", -- Line 1   Column 3535   Coefficient 70.96777344
   "010001101111100010", -- Line 1   Column 3536   Coefficient 70.97070313
   "010001101111100100", -- Line 1   Column 3537   Coefficient 70.97265625
   "010001101111100111", -- Line 1   Column 3538   Coefficient 70.97558594
   "010001101111101001", -- Line 1   Column 3539   Coefficient 70.97753906
   "010001101111101100", -- Line 1   Column 3540   Coefficient 70.98046875
   "010001101111101110", -- Line 1   Column 3541   Coefficient 70.98242188
   "010001101111110001", -- Line 1   Column 3542   Coefficient 70.98535156
   "010001101111110011", -- Line 1   Column 3543   Coefficient 70.98730469
   "010001101111110110", -- Line 1   Column 3544   Coefficient 70.99023438
   "010001101111111000", -- Line 1   Column 3545   Coefficient 70.99218750
   "010001101111111011", -- Line 1   Column 3546   Coefficient 70.99511719
   "010001101111111101", -- Line 1   Column 3547   Coefficient 70.99707031
   "010001110000000000", -- Line 1   Column 3548   Coefficient 71.00000000
   "010001110000000010", -- Line 1   Column 3549   Coefficient 71.00195313
   "010001110000000101", -- Line 1   Column 3550   Coefficient 71.00488281
   "010001110000000111", -- Line 1   Column 3551   Coefficient 71.00683594
   "010001110000001010", -- Line 1   Column 3552   Coefficient 71.00976563
   "010001110000001100", -- Line 1   Column 3553   Coefficient 71.01171875
   "010001110000001111", -- Line 1   Column 3554   Coefficient 71.01464844
   "010001110000010001", -- Line 1   Column 3555   Coefficient 71.01660156
   "010001110000010100", -- Line 1   Column 3556   Coefficient 71.01953125
   "010001110000010110", -- Line 1   Column 3557   Coefficient 71.02148438
   "010001110000011001", -- Line 1   Column 3558   Coefficient 71.02441406
   "010001110000011011", -- Line 1   Column 3559   Coefficient 71.02636719
   "010001110000011110", -- Line 1   Column 3560   Coefficient 71.02929688
   "010001110000100000", -- Line 1   Column 3561   Coefficient 71.03125000
   "010001110000100011", -- Line 1   Column 3562   Coefficient 71.03417969
   "010001110000100101", -- Line 1   Column 3563   Coefficient 71.03613281
   "010001110000101000", -- Line 1   Column 3564   Coefficient 71.03906250
   "010001110000101010", -- Line 1   Column 3565   Coefficient 71.04101563
   "010001110000101101", -- Line 1   Column 3566   Coefficient 71.04394531
   "010001110000101111", -- Line 1   Column 3567   Coefficient 71.04589844
   "010001110000110010", -- Line 1   Column 3568   Coefficient 71.04882813
   "010001110000110100", -- Line 1   Column 3569   Coefficient 71.05078125
   "010001110000110111", -- Line 1   Column 3570   Coefficient 71.05371094
   "010001110000111001", -- Line 1   Column 3571   Coefficient 71.05566406
   "010001110000111100", -- Line 1   Column 3572   Coefficient 71.05859375
   "010001110000111110", -- Line 1   Column 3573   Coefficient 71.06054688
   "010001110001000001", -- Line 1   Column 3574   Coefficient 71.06347656
   "010001110001000011", -- Line 1   Column 3575   Coefficient 71.06542969
   "010001110001000110", -- Line 1   Column 3576   Coefficient 71.06835938
   "010001110001001000", -- Line 1   Column 3577   Coefficient 71.07031250
   "010001110001001011", -- Line 1   Column 3578   Coefficient 71.07324219
   "010001110001001101", -- Line 1   Column 3579   Coefficient 71.07519531
   "010001110001010000", -- Line 1   Column 3580   Coefficient 71.07812500
   "010001110001010010", -- Line 1   Column 3581   Coefficient 71.08007813
   "010001110001010100", -- Line 1   Column 3582   Coefficient 71.08203125
   "010001110001010111", -- Line 1   Column 3583   Coefficient 71.08496094
   "010001110001011001", -- Line 1   Column 3584   Coefficient 71.08691406
   "010001110001011100", -- Line 1   Column 3585   Coefficient 71.08984375
   "010001110001011110", -- Line 1   Column 3586   Coefficient 71.09179688
   "010001110001100001", -- Line 1   Column 3587   Coefficient 71.09472656
   "010001110001100011", -- Line 1   Column 3588   Coefficient 71.09667969
   "010001110001100110", -- Line 1   Column 3589   Coefficient 71.09960938
   "010001110001101000", -- Line 1   Column 3590   Coefficient 71.10156250
   "010001110001101011", -- Line 1   Column 3591   Coefficient 71.10449219
   "010001110001101101", -- Line 1   Column 3592   Coefficient 71.10644531
   "010001110001110000", -- Line 1   Column 3593   Coefficient 71.10937500
   "010001110001110010", -- Line 1   Column 3594   Coefficient 71.11132813
   "010001110001110101", -- Line 1   Column 3595   Coefficient 71.11425781
   "010001110001110111", -- Line 1   Column 3596   Coefficient 71.11621094
   "010001110001111010", -- Line 1   Column 3597   Coefficient 71.11914063
   "010001110001111100", -- Line 1   Column 3598   Coefficient 71.12109375
   "010001110001111111", -- Line 1   Column 3599   Coefficient 71.12402344
   "010001110010000001", -- Line 1   Column 3600   Coefficient 71.12597656
   "010001110010000100", -- Line 1   Column 3601   Coefficient 71.12890625
   "010001110010000110", -- Line 1   Column 3602   Coefficient 71.13085938
   "010001110010001000", -- Line 1   Column 3603   Coefficient 71.13281250
   "010001110010001011", -- Line 1   Column 3604   Coefficient 71.13574219
   "010001110010001101", -- Line 1   Column 3605   Coefficient 71.13769531
   "010001110010010000", -- Line 1   Column 3606   Coefficient 71.14062500
   "010001110010010010", -- Line 1   Column 3607   Coefficient 71.14257813
   "010001110010010101", -- Line 1   Column 3608   Coefficient 71.14550781
   "010001110010010111", -- Line 1   Column 3609   Coefficient 71.14746094
   "010001110010011010", -- Line 1   Column 3610   Coefficient 71.15039063
   "010001110010011100", -- Line 1   Column 3611   Coefficient 71.15234375
   "010001110010011111", -- Line 1   Column 3612   Coefficient 71.15527344
   "010001110010100001", -- Line 1   Column 3613   Coefficient 71.15722656
   "010001110010100100", -- Line 1   Column 3614   Coefficient 71.16015625
   "010001110010100110", -- Line 1   Column 3615   Coefficient 71.16210938
   "010001110010101001", -- Line 1   Column 3616   Coefficient 71.16503906
   "010001110010101011", -- Line 1   Column 3617   Coefficient 71.16699219
   "010001110010101101", -- Line 1   Column 3618   Coefficient 71.16894531
   "010001110010110000", -- Line 1   Column 3619   Coefficient 71.17187500
   "010001110010110010", -- Line 1   Column 3620   Coefficient 71.17382813
   "010001110010110101", -- Line 1   Column 3621   Coefficient 71.17675781
   "010001110010110111", -- Line 1   Column 3622   Coefficient 71.17871094
   "010001110010111010", -- Line 1   Column 3623   Coefficient 71.18164063
   "010001110010111100", -- Line 1   Column 3624   Coefficient 71.18359375
   "010001110010111111", -- Line 1   Column 3625   Coefficient 71.18652344
   "010001110011000001", -- Line 1   Column 3626   Coefficient 71.18847656
   "010001110011000100", -- Line 1   Column 3627   Coefficient 71.19140625
   "010001110011000110", -- Line 1   Column 3628   Coefficient 71.19335938
   "010001110011001000", -- Line 1   Column 3629   Coefficient 71.19531250
   "010001110011001011", -- Line 1   Column 3630   Coefficient 71.19824219
   "010001110011001101", -- Line 1   Column 3631   Coefficient 71.20019531
   "010001110011010000", -- Line 1   Column 3632   Coefficient 71.20312500
   "010001110011010010", -- Line 1   Column 3633   Coefficient 71.20507813
   "010001110011010101", -- Line 1   Column 3634   Coefficient 71.20800781
   "010001110011010111", -- Line 1   Column 3635   Coefficient 71.20996094
   "010001110011011010", -- Line 1   Column 3636   Coefficient 71.21289063
   "010001110011011100", -- Line 1   Column 3637   Coefficient 71.21484375
   "010001110011011110", -- Line 1   Column 3638   Coefficient 71.21679688
   "010001110011100001", -- Line 1   Column 3639   Coefficient 71.21972656
   "010001110011100011", -- Line 1   Column 3640   Coefficient 71.22167969
   "010001110011100110", -- Line 1   Column 3641   Coefficient 71.22460938
   "010001110011101000", -- Line 1   Column 3642   Coefficient 71.22656250
   "010001110011101011", -- Line 1   Column 3643   Coefficient 71.22949219
   "010001110011101101", -- Line 1   Column 3644   Coefficient 71.23144531
   "010001110011110000", -- Line 1   Column 3645   Coefficient 71.23437500
   "010001110011110010", -- Line 1   Column 3646   Coefficient 71.23632813
   "010001110011110100", -- Line 1   Column 3647   Coefficient 71.23828125
   "010001110011110111", -- Line 1   Column 3648   Coefficient 71.24121094
   "010001110011111001", -- Line 1   Column 3649   Coefficient 71.24316406
   "010001110011111100", -- Line 1   Column 3650   Coefficient 71.24609375
   "010001110011111110", -- Line 1   Column 3651   Coefficient 71.24804688
   "010001110100000001", -- Line 1   Column 3652   Coefficient 71.25097656
   "010001110100000011", -- Line 1   Column 3653   Coefficient 71.25292969
   "010001110100000101", -- Line 1   Column 3654   Coefficient 71.25488281
   "010001110100001000", -- Line 1   Column 3655   Coefficient 71.25781250
   "010001110100001010", -- Line 1   Column 3656   Coefficient 71.25976563
   "010001110100001101", -- Line 1   Column 3657   Coefficient 71.26269531
   "010001110100001111", -- Line 1   Column 3658   Coefficient 71.26464844
   "010001110100010010", -- Line 1   Column 3659   Coefficient 71.26757813
   "010001110100010100", -- Line 1   Column 3660   Coefficient 71.26953125
   "010001110100010111", -- Line 1   Column 3661   Coefficient 71.27246094
   "010001110100011001", -- Line 1   Column 3662   Coefficient 71.27441406
   "010001110100011011", -- Line 1   Column 3663   Coefficient 71.27636719
   "010001110100011110", -- Line 1   Column 3664   Coefficient 71.27929688
   "010001110100100000", -- Line 1   Column 3665   Coefficient 71.28125000
   "010001110100100011", -- Line 1   Column 3666   Coefficient 71.28417969
   "010001110100100101", -- Line 1   Column 3667   Coefficient 71.28613281
   "010001110100101000", -- Line 1   Column 3668   Coefficient 71.28906250
   "010001110100101010", -- Line 1   Column 3669   Coefficient 71.29101563
   "010001110100101100", -- Line 1   Column 3670   Coefficient 71.29296875
   "010001110100101111", -- Line 1   Column 3671   Coefficient 71.29589844
   "010001110100110001", -- Line 1   Column 3672   Coefficient 71.29785156
   "010001110100110100", -- Line 1   Column 3673   Coefficient 71.30078125
   "010001110100110110", -- Line 1   Column 3674   Coefficient 71.30273438
   "010001110100111000", -- Line 1   Column 3675   Coefficient 71.30468750
   "010001110100111011", -- Line 1   Column 3676   Coefficient 71.30761719
   "010001110100111101", -- Line 1   Column 3677   Coefficient 71.30957031
   "010001110101000000", -- Line 1   Column 3678   Coefficient 71.31250000
   "010001110101000010", -- Line 1   Column 3679   Coefficient 71.31445313
   "010001110101000101", -- Line 1   Column 3680   Coefficient 71.31738281
   "010001110101000111", -- Line 1   Column 3681   Coefficient 71.31933594
   "010001110101001001", -- Line 1   Column 3682   Coefficient 71.32128906
   "010001110101001100", -- Line 1   Column 3683   Coefficient 71.32421875
   "010001110101001110", -- Line 1   Column 3684   Coefficient 71.32617188
   "010001110101010001", -- Line 1   Column 3685   Coefficient 71.32910156
   "010001110101010011", -- Line 1   Column 3686   Coefficient 71.33105469
   "010001110101010101", -- Line 1   Column 3687   Coefficient 71.33300781
   "010001110101011000", -- Line 1   Column 3688   Coefficient 71.33593750
   "010001110101011010", -- Line 1   Column 3689   Coefficient 71.33789063
   "010001110101011101", -- Line 1   Column 3690   Coefficient 71.34082031
   "010001110101011111", -- Line 1   Column 3691   Coefficient 71.34277344
   "010001110101100010", -- Line 1   Column 3692   Coefficient 71.34570313
   "010001110101100100", -- Line 1   Column 3693   Coefficient 71.34765625
   "010001110101100110", -- Line 1   Column 3694   Coefficient 71.34960938
   "010001110101101001", -- Line 1   Column 3695   Coefficient 71.35253906
   "010001110101101011", -- Line 1   Column 3696   Coefficient 71.35449219
   "010001110101101110", -- Line 1   Column 3697   Coefficient 71.35742188
   "010001110101110000", -- Line 1   Column 3698   Coefficient 71.35937500
   "010001110101110010", -- Line 1   Column 3699   Coefficient 71.36132813
   "010001110101110101", -- Line 1   Column 3700   Coefficient 71.36425781
   "010001110101110111", -- Line 1   Column 3701   Coefficient 71.36621094
   "010001110101111010", -- Line 1   Column 3702   Coefficient 71.36914063
   "010001110101111100", -- Line 1   Column 3703   Coefficient 71.37109375
   "010001110101111110", -- Line 1   Column 3704   Coefficient 71.37304688
   "010001110110000001", -- Line 1   Column 3705   Coefficient 71.37597656
   "010001110110000011", -- Line 1   Column 3706   Coefficient 71.37792969
   "010001110110000110", -- Line 1   Column 3707   Coefficient 71.38085938
   "010001110110001000", -- Line 1   Column 3708   Coefficient 71.38281250
   "010001110110001010", -- Line 1   Column 3709   Coefficient 71.38476563
   "010001110110001101", -- Line 1   Column 3710   Coefficient 71.38769531
   "010001110110001111", -- Line 1   Column 3711   Coefficient 71.38964844
   "010001110110010010", -- Line 1   Column 3712   Coefficient 71.39257813
   "010001110110010100", -- Line 1   Column 3713   Coefficient 71.39453125
   "010001110110010110", -- Line 1   Column 3714   Coefficient 71.39648438
   "010001110110011001", -- Line 1   Column 3715   Coefficient 71.39941406
   "010001110110011011", -- Line 1   Column 3716   Coefficient 71.40136719
   "010001110110011110", -- Line 1   Column 3717   Coefficient 71.40429688
   "010001110110100000", -- Line 1   Column 3718   Coefficient 71.40625000
   "010001110110100010", -- Line 1   Column 3719   Coefficient 71.40820313
   "010001110110100101", -- Line 1   Column 3720   Coefficient 71.41113281
   "010001110110100111", -- Line 1   Column 3721   Coefficient 71.41308594
   "010001110110101010", -- Line 1   Column 3722   Coefficient 71.41601563
   "010001110110101100", -- Line 1   Column 3723   Coefficient 71.41796875
   "010001110110101110", -- Line 1   Column 3724   Coefficient 71.41992188
   "010001110110110001", -- Line 1   Column 3725   Coefficient 71.42285156
   "010001110110110011", -- Line 1   Column 3726   Coefficient 71.42480469
   "010001110110110101", -- Line 1   Column 3727   Coefficient 71.42675781
   "010001110110111000", -- Line 1   Column 3728   Coefficient 71.42968750
   "010001110110111010", -- Line 1   Column 3729   Coefficient 71.43164063
   "010001110110111101", -- Line 1   Column 3730   Coefficient 71.43457031
   "010001110110111111", -- Line 1   Column 3731   Coefficient 71.43652344
   "010001110111000001", -- Line 1   Column 3732   Coefficient 71.43847656
   "010001110111000100", -- Line 1   Column 3733   Coefficient 71.44140625
   "010001110111000110", -- Line 1   Column 3734   Coefficient 71.44335938
   "010001110111001001", -- Line 1   Column 3735   Coefficient 71.44628906
   "010001110111001011", -- Line 1   Column 3736   Coefficient 71.44824219
   "010001110111001101", -- Line 1   Column 3737   Coefficient 71.45019531
   "010001110111010000", -- Line 1   Column 3738   Coefficient 71.45312500
   "010001110111010010", -- Line 1   Column 3739   Coefficient 71.45507813
   "010001110111010100", -- Line 1   Column 3740   Coefficient 71.45703125
   "010001110111010111", -- Line 1   Column 3741   Coefficient 71.45996094
   "010001110111011001", -- Line 1   Column 3742   Coefficient 71.46191406
   "010001110111011100", -- Line 1   Column 3743   Coefficient 71.46484375
   "010001110111011110", -- Line 1   Column 3744   Coefficient 71.46679688
   "010001110111100000", -- Line 1   Column 3745   Coefficient 71.46875000
   "010001110111100011", -- Line 1   Column 3746   Coefficient 71.47167969
   "010001110111100101", -- Line 1   Column 3747   Coefficient 71.47363281
   "010001110111100111", -- Line 1   Column 3748   Coefficient 71.47558594
   "010001110111101010", -- Line 1   Column 3749   Coefficient 71.47851563
   "010001110111101100", -- Line 1   Column 3750   Coefficient 71.48046875
   "010001110111101111", -- Line 1   Column 3751   Coefficient 71.48339844
   "010001110111110001", -- Line 1   Column 3752   Coefficient 71.48535156
   "010001110111110011", -- Line 1   Column 3753   Coefficient 71.48730469
   "010001110111110110", -- Line 1   Column 3754   Coefficient 71.49023438
   "010001110111111000", -- Line 1   Column 3755   Coefficient 71.49218750
   "010001110111111010", -- Line 1   Column 3756   Coefficient 71.49414063
   "010001110111111101", -- Line 1   Column 3757   Coefficient 71.49707031
   "010001110111111111", -- Line 1   Column 3758   Coefficient 71.49902344
   "010001111000000001", -- Line 1   Column 3759   Coefficient 71.50097656
   "010001111000000100", -- Line 1   Column 3760   Coefficient 71.50390625
   "010001111000000110", -- Line 1   Column 3761   Coefficient 71.50585938
   "010001111000001001", -- Line 1   Column 3762   Coefficient 71.50878906
   "010001111000001011", -- Line 1   Column 3763   Coefficient 71.51074219
   "010001111000001101", -- Line 1   Column 3764   Coefficient 71.51269531
   "010001111000010000", -- Line 1   Column 3765   Coefficient 71.51562500
   "010001111000010010", -- Line 1   Column 3766   Coefficient 71.51757813
   "010001111000010100", -- Line 1   Column 3767   Coefficient 71.51953125
   "010001111000010111", -- Line 1   Column 3768   Coefficient 71.52246094
   "010001111000011001", -- Line 1   Column 3769   Coefficient 71.52441406
   "010001111000011011", -- Line 1   Column 3770   Coefficient 71.52636719
   "010001111000011110", -- Line 1   Column 3771   Coefficient 71.52929688
   "010001111000100000", -- Line 1   Column 3772   Coefficient 71.53125000
   "010001111000100011", -- Line 1   Column 3773   Coefficient 71.53417969
   "010001111000100101", -- Line 1   Column 3774   Coefficient 71.53613281
   "010001111000100111", -- Line 1   Column 3775   Coefficient 71.53808594
   "010001111000101010", -- Line 1   Column 3776   Coefficient 71.54101563
   "010001111000101100", -- Line 1   Column 3777   Coefficient 71.54296875
   "010001111000101110", -- Line 1   Column 3778   Coefficient 71.54492188
   "010001111000110001", -- Line 1   Column 3779   Coefficient 71.54785156
   "010001111000110011", -- Line 1   Column 3780   Coefficient 71.54980469
   "010001111000110101", -- Line 1   Column 3781   Coefficient 71.55175781
   "010001111000111000", -- Line 1   Column 3782   Coefficient 71.55468750
   "010001111000111010", -- Line 1   Column 3783   Coefficient 71.55664063
   "010001111000111100", -- Line 1   Column 3784   Coefficient 71.55859375
   "010001111000111111", -- Line 1   Column 3785   Coefficient 71.56152344
   "010001111001000001", -- Line 1   Column 3786   Coefficient 71.56347656
   "010001111001000011", -- Line 1   Column 3787   Coefficient 71.56542969
   "010001111001000110", -- Line 1   Column 3788   Coefficient 71.56835938
   "010001111001001000", -- Line 1   Column 3789   Coefficient 71.57031250
   "010001111001001011", -- Line 1   Column 3790   Coefficient 71.57324219
   "010001111001001101", -- Line 1   Column 3791   Coefficient 71.57519531
   "010001111001001111", -- Line 1   Column 3792   Coefficient 71.57714844
   "010001111001010010", -- Line 1   Column 3793   Coefficient 71.58007813
   "010001111001010100", -- Line 1   Column 3794   Coefficient 71.58203125
   "010001111001010110", -- Line 1   Column 3795   Coefficient 71.58398438
   "010001111001011001", -- Line 1   Column 3796   Coefficient 71.58691406
   "010001111001011011", -- Line 1   Column 3797   Coefficient 71.58886719
   "010001111001011101", -- Line 1   Column 3798   Coefficient 71.59082031
   "010001111001100000", -- Line 1   Column 3799   Coefficient 71.59375000
   "010001111001100010", -- Line 1   Column 3800   Coefficient 71.59570313
   "010001111001100100", -- Line 1   Column 3801   Coefficient 71.59765625
   "010001111001100111", -- Line 1   Column 3802   Coefficient 71.60058594
   "010001111001101001", -- Line 1   Column 3803   Coefficient 71.60253906
   "010001111001101011", -- Line 1   Column 3804   Coefficient 71.60449219
   "010001111001101110", -- Line 1   Column 3805   Coefficient 71.60742188
   "010001111001110000", -- Line 1   Column 3806   Coefficient 71.60937500
   "010001111001110010", -- Line 1   Column 3807   Coefficient 71.61132813
   "010001111001110101", -- Line 1   Column 3808   Coefficient 71.61425781
   "010001111001110111", -- Line 1   Column 3809   Coefficient 71.61621094
   "010001111001111001", -- Line 1   Column 3810   Coefficient 71.61816406
   "010001111001111100", -- Line 1   Column 3811   Coefficient 71.62109375
   "010001111001111110", -- Line 1   Column 3812   Coefficient 71.62304688
   "010001111010000000", -- Line 1   Column 3813   Coefficient 71.62500000
   "010001111010000011", -- Line 1   Column 3814   Coefficient 71.62792969
   "010001111010000101", -- Line 1   Column 3815   Coefficient 71.62988281
   "010001111010000111", -- Line 1   Column 3816   Coefficient 71.63183594
   "010001111010001010", -- Line 1   Column 3817   Coefficient 71.63476563
   "010001111010001100", -- Line 1   Column 3818   Coefficient 71.63671875
   "010001111010001110", -- Line 1   Column 3819   Coefficient 71.63867188
   "010001111010010001", -- Line 1   Column 3820   Coefficient 71.64160156
   "010001111010010011", -- Line 1   Column 3821   Coefficient 71.64355469
   "010001111010010101", -- Line 1   Column 3822   Coefficient 71.64550781
   "010001111010011000", -- Line 1   Column 3823   Coefficient 71.64843750
   "010001111010011010", -- Line 1   Column 3824   Coefficient 71.65039063
   "010001111010011100", -- Line 1   Column 3825   Coefficient 71.65234375
   "010001111010011111", -- Line 1   Column 3826   Coefficient 71.65527344
   "010001111010100001", -- Line 1   Column 3827   Coefficient 71.65722656
   "010001111010100011", -- Line 1   Column 3828   Coefficient 71.65917969
   "010001111010100110", -- Line 1   Column 3829   Coefficient 71.66210938
   "010001111010101000", -- Line 1   Column 3830   Coefficient 71.66406250
   "010001111010101010", -- Line 1   Column 3831   Coefficient 71.66601563
   "010001111010101101", -- Line 1   Column 3832   Coefficient 71.66894531
   "010001111010101111", -- Line 1   Column 3833   Coefficient 71.67089844
   "010001111010110001", -- Line 1   Column 3834   Coefficient 71.67285156
   "010001111010110100", -- Line 1   Column 3835   Coefficient 71.67578125
   "010001111010110110", -- Line 1   Column 3836   Coefficient 71.67773438
   "010001111010111000", -- Line 1   Column 3837   Coefficient 71.67968750
   "010001111010111010", -- Line 1   Column 3838   Coefficient 71.68164063
   "010001111010111101", -- Line 1   Column 3839   Coefficient 71.68457031
   "010001111010111111", -- Line 1   Column 3840   Coefficient 71.68652344
   "010001111011000001", -- Line 1   Column 3841   Coefficient 71.68847656
   "010001111011000100", -- Line 1   Column 3842   Coefficient 71.69140625
   "010001111011000110", -- Line 1   Column 3843   Coefficient 71.69335938
   "010001111011001000", -- Line 1   Column 3844   Coefficient 71.69531250
   "010001111011001011", -- Line 1   Column 3845   Coefficient 71.69824219
   "010001111011001101", -- Line 1   Column 3846   Coefficient 71.70019531
   "010001111011001111", -- Line 1   Column 3847   Coefficient 71.70214844
   "010001111011010010", -- Line 1   Column 3848   Coefficient 71.70507813
   "010001111011010100", -- Line 1   Column 3849   Coefficient 71.70703125
   "010001111011010110", -- Line 1   Column 3850   Coefficient 71.70898438
   "010001111011011001", -- Line 1   Column 3851   Coefficient 71.71191406
   "010001111011011011", -- Line 1   Column 3852   Coefficient 71.71386719
   "010001111011011101", -- Line 1   Column 3853   Coefficient 71.71582031
   "010001111011011111", -- Line 1   Column 3854   Coefficient 71.71777344
   "010001111011100010", -- Line 1   Column 3855   Coefficient 71.72070313
   "010001111011100100", -- Line 1   Column 3856   Coefficient 71.72265625
   "010001111011100110", -- Line 1   Column 3857   Coefficient 71.72460938
   "010001111011101001", -- Line 1   Column 3858   Coefficient 71.72753906
   "010001111011101011", -- Line 1   Column 3859   Coefficient 71.72949219
   "010001111011101101", -- Line 1   Column 3860   Coefficient 71.73144531
   "010001111011110000", -- Line 1   Column 3861   Coefficient 71.73437500
   "010001111011110010", -- Line 1   Column 3862   Coefficient 71.73632813
   "010001111011110100", -- Line 1   Column 3863   Coefficient 71.73828125
   "010001111011110111", -- Line 1   Column 3864   Coefficient 71.74121094
   "010001111011111001", -- Line 1   Column 3865   Coefficient 71.74316406
   "010001111011111011", -- Line 1   Column 3866   Coefficient 71.74511719
   "010001111011111101", -- Line 1   Column 3867   Coefficient 71.74707031
   "010001111100000000", -- Line 1   Column 3868   Coefficient 71.75000000
   "010001111100000010", -- Line 1   Column 3869   Coefficient 71.75195313
   "010001111100000100", -- Line 1   Column 3870   Coefficient 71.75390625
   "010001111100000111", -- Line 1   Column 3871   Coefficient 71.75683594
   "010001111100001001", -- Line 1   Column 3872   Coefficient 71.75878906
   "010001111100001011", -- Line 1   Column 3873   Coefficient 71.76074219
   "010001111100001110", -- Line 1   Column 3874   Coefficient 71.76367188
   "010001111100010000", -- Line 1   Column 3875   Coefficient 71.76562500
   "010001111100010010", -- Line 1   Column 3876   Coefficient 71.76757813
   "010001111100010100", -- Line 1   Column 3877   Coefficient 71.76953125
   "010001111100010111", -- Line 1   Column 3878   Coefficient 71.77246094
   "010001111100011001", -- Line 1   Column 3879   Coefficient 71.77441406
   "010001111100011011", -- Line 1   Column 3880   Coefficient 71.77636719
   "010001111100011110", -- Line 1   Column 3881   Coefficient 71.77929688
   "010001111100100000", -- Line 1   Column 3882   Coefficient 71.78125000
   "010001111100100010", -- Line 1   Column 3883   Coefficient 71.78320313
   "010001111100100100", -- Line 1   Column 3884   Coefficient 71.78515625
   "010001111100100111", -- Line 1   Column 3885   Coefficient 71.78808594
   "010001111100101001", -- Line 1   Column 3886   Coefficient 71.79003906
   "010001111100101011", -- Line 1   Column 3887   Coefficient 71.79199219
   "010001111100101110", -- Line 1   Column 3888   Coefficient 71.79492188
   "010001111100110000", -- Line 1   Column 3889   Coefficient 71.79687500
   "010001111100110010", -- Line 1   Column 3890   Coefficient 71.79882813
   "010001111100110100", -- Line 1   Column 3891   Coefficient 71.80078125
   "010001111100110111", -- Line 1   Column 3892   Coefficient 71.80371094
   "010001111100111001", -- Line 1   Column 3893   Coefficient 71.80566406
   "010001111100111011", -- Line 1   Column 3894   Coefficient 71.80761719
   "010001111100111110", -- Line 1   Column 3895   Coefficient 71.81054688
   "010001111101000000", -- Line 1   Column 3896   Coefficient 71.81250000
   "010001111101000010", -- Line 1   Column 3897   Coefficient 71.81445313
   "010001111101000100", -- Line 1   Column 3898   Coefficient 71.81640625
   "010001111101000111", -- Line 1   Column 3899   Coefficient 71.81933594
   "010001111101001001", -- Line 1   Column 3900   Coefficient 71.82128906
   "010001111101001011", -- Line 1   Column 3901   Coefficient 71.82324219
   "010001111101001110", -- Line 1   Column 3902   Coefficient 71.82617188
   "010001111101010000", -- Line 1   Column 3903   Coefficient 71.82812500
   "010001111101010010", -- Line 1   Column 3904   Coefficient 71.83007813
   "010001111101010100", -- Line 1   Column 3905   Coefficient 71.83203125
   "010001111101010111", -- Line 1   Column 3906   Coefficient 71.83496094
   "010001111101011001", -- Line 1   Column 3907   Coefficient 71.83691406
   "010001111101011011", -- Line 1   Column 3908   Coefficient 71.83886719
   "010001111101011110", -- Line 1   Column 3909   Coefficient 71.84179688
   "010001111101100000", -- Line 1   Column 3910   Coefficient 71.84375000
   "010001111101100010", -- Line 1   Column 3911   Coefficient 71.84570313
   "010001111101100100", -- Line 1   Column 3912   Coefficient 71.84765625
   "010001111101100111", -- Line 1   Column 3913   Coefficient 71.85058594
   "010001111101101001", -- Line 1   Column 3914   Coefficient 71.85253906
   "010001111101101011", -- Line 1   Column 3915   Coefficient 71.85449219
   "010001111101101101", -- Line 1   Column 3916   Coefficient 71.85644531
   "010001111101110000", -- Line 1   Column 3917   Coefficient 71.85937500
   "010001111101110010", -- Line 1   Column 3918   Coefficient 71.86132813
   "010001111101110100", -- Line 1   Column 3919   Coefficient 71.86328125
   "010001111101110110", -- Line 1   Column 3920   Coefficient 71.86523438
   "010001111101111001", -- Line 1   Column 3921   Coefficient 71.86816406
   "010001111101111011", -- Line 1   Column 3922   Coefficient 71.87011719
   "010001111101111101", -- Line 1   Column 3923   Coefficient 71.87207031
   "010001111110000000", -- Line 1   Column 3924   Coefficient 71.87500000
   "010001111110000010", -- Line 1   Column 3925   Coefficient 71.87695313
   "010001111110000100", -- Line 1   Column 3926   Coefficient 71.87890625
   "010001111110000110", -- Line 1   Column 3927   Coefficient 71.88085938
   "010001111110001001", -- Line 1   Column 3928   Coefficient 71.88378906
   "010001111110001011", -- Line 1   Column 3929   Coefficient 71.88574219
   "010001111110001101", -- Line 1   Column 3930   Coefficient 71.88769531
   "010001111110001111", -- Line 1   Column 3931   Coefficient 71.88964844
   "010001111110010010", -- Line 1   Column 3932   Coefficient 71.89257813
   "010001111110010100", -- Line 1   Column 3933   Coefficient 71.89453125
   "010001111110010110", -- Line 1   Column 3934   Coefficient 71.89648438
   "010001111110011000", -- Line 1   Column 3935   Coefficient 71.89843750
   "010001111110011011", -- Line 1   Column 3936   Coefficient 71.90136719
   "010001111110011101", -- Line 1   Column 3937   Coefficient 71.90332031
   "010001111110011111", -- Line 1   Column 3938   Coefficient 71.90527344
   "010001111110100010", -- Line 1   Column 3939   Coefficient 71.90820313
   "010001111110100100", -- Line 1   Column 3940   Coefficient 71.91015625
   "010001111110100110", -- Line 1   Column 3941   Coefficient 71.91210938
   "010001111110101000", -- Line 1   Column 3942   Coefficient 71.91406250
   "010001111110101011", -- Line 1   Column 3943   Coefficient 71.91699219
   "010001111110101101", -- Line 1   Column 3944   Coefficient 71.91894531
   "010001111110101111", -- Line 1   Column 3945   Coefficient 71.92089844
   "010001111110110001", -- Line 1   Column 3946   Coefficient 71.92285156
   "010001111110110100", -- Line 1   Column 3947   Coefficient 71.92578125
   "010001111110110110", -- Line 1   Column 3948   Coefficient 71.92773438
   "010001111110111000", -- Line 1   Column 3949   Coefficient 71.92968750
   "010001111110111010", -- Line 1   Column 3950   Coefficient 71.93164063
   "010001111110111101", -- Line 1   Column 3951   Coefficient 71.93457031
   "010001111110111111", -- Line 1   Column 3952   Coefficient 71.93652344
   "010001111111000001", -- Line 1   Column 3953   Coefficient 71.93847656
   "010001111111000011", -- Line 1   Column 3954   Coefficient 71.94042969
   "010001111111000110", -- Line 1   Column 3955   Coefficient 71.94335938
   "010001111111001000", -- Line 1   Column 3956   Coefficient 71.94531250
   "010001111111001010", -- Line 1   Column 3957   Coefficient 71.94726563
   "010001111111001100", -- Line 1   Column 3958   Coefficient 71.94921875
   "010001111111001111", -- Line 1   Column 3959   Coefficient 71.95214844
   "010001111111010001", -- Line 1   Column 3960   Coefficient 71.95410156
   "010001111111010011", -- Line 1   Column 3961   Coefficient 71.95605469
   "010001111111010101", -- Line 1   Column 3962   Coefficient 71.95800781
   "010001111111011000", -- Line 1   Column 3963   Coefficient 71.96093750
   "010001111111011010", -- Line 1   Column 3964   Coefficient 71.96289063
   "010001111111011100", -- Line 1   Column 3965   Coefficient 71.96484375
   "010001111111011110", -- Line 1   Column 3966   Coefficient 71.96679688
   "010001111111100001", -- Line 1   Column 3967   Coefficient 71.96972656
   "010001111111100011", -- Line 1   Column 3968   Coefficient 71.97167969
   "010001111111100101", -- Line 1   Column 3969   Coefficient 71.97363281
   "010001111111100111", -- Line 1   Column 3970   Coefficient 71.97558594
   "010001111111101001", -- Line 1   Column 3971   Coefficient 71.97753906
   "010001111111101100", -- Line 1   Column 3972   Coefficient 71.98046875
   "010001111111101110", -- Line 1   Column 3973   Coefficient 71.98242188
   "010001111111110000", -- Line 1   Column 3974   Coefficient 71.98437500
   "010001111111110010", -- Line 1   Column 3975   Coefficient 71.98632813
   "010001111111110101", -- Line 1   Column 3976   Coefficient 71.98925781
   "010001111111110111", -- Line 1   Column 3977   Coefficient 71.99121094
   "010001111111111001", -- Line 1   Column 3978   Coefficient 71.99316406
   "010001111111111011", -- Line 1   Column 3979   Coefficient 71.99511719
   "010001111111111110", -- Line 1   Column 3980   Coefficient 71.99804688
   "010010000000000000", -- Line 1   Column 3981   Coefficient 72.00000000
   "010010000000000010", -- Line 1   Column 3982   Coefficient 72.00195313
   "010010000000000100", -- Line 1   Column 3983   Coefficient 72.00390625
   "010010000000000111", -- Line 1   Column 3984   Coefficient 72.00683594
   "010010000000001001", -- Line 1   Column 3985   Coefficient 72.00878906
   "010010000000001011", -- Line 1   Column 3986   Coefficient 72.01074219
   "010010000000001101", -- Line 1   Column 3987   Coefficient 72.01269531
   "010010000000001111", -- Line 1   Column 3988   Coefficient 72.01464844
   "010010000000010010", -- Line 1   Column 3989   Coefficient 72.01757813
   "010010000000010100", -- Line 1   Column 3990   Coefficient 72.01953125
   "010010000000010110", -- Line 1   Column 3991   Coefficient 72.02148438
   "010010000000011000", -- Line 1   Column 3992   Coefficient 72.02343750
   "010010000000011011", -- Line 1   Column 3993   Coefficient 72.02636719
   "010010000000011101", -- Line 1   Column 3994   Coefficient 72.02832031
   "010010000000011111", -- Line 1   Column 3995   Coefficient 72.03027344
   "010010000000100001", -- Line 1   Column 3996   Coefficient 72.03222656
   "010010000000100100", -- Line 1   Column 3997   Coefficient 72.03515625
   "010010000000100110", -- Line 1   Column 3998   Coefficient 72.03710938
   "010010000000101000", -- Line 1   Column 3999   Coefficient 72.03906250
   "010010000000101010", -- Line 1   Column 4000   Coefficient 72.04101563
   "010010000000101100", -- Line 1   Column 4001   Coefficient 72.04296875
   "010010000000101111", -- Line 1   Column 4002   Coefficient 72.04589844
   "010010000000110001", -- Line 1   Column 4003   Coefficient 72.04785156
   "010010000000110011", -- Line 1   Column 4004   Coefficient 72.04980469
   "010010000000110101", -- Line 1   Column 4005   Coefficient 72.05175781
   "010010000000111000", -- Line 1   Column 4006   Coefficient 72.05468750
   "010010000000111010", -- Line 1   Column 4007   Coefficient 72.05664063
   "010010000000111100", -- Line 1   Column 4008   Coefficient 72.05859375
   "010010000000111110", -- Line 1   Column 4009   Coefficient 72.06054688
   "010010000001000000", -- Line 1   Column 4010   Coefficient 72.06250000
   "010010000001000011", -- Line 1   Column 4011   Coefficient 72.06542969
   "010010000001000101", -- Line 1   Column 4012   Coefficient 72.06738281
   "010010000001000111", -- Line 1   Column 4013   Coefficient 72.06933594
   "010010000001001001", -- Line 1   Column 4014   Coefficient 72.07128906
   "010010000001001011", -- Line 1   Column 4015   Coefficient 72.07324219
   "010010000001001110", -- Line 1   Column 4016   Coefficient 72.07617188
   "010010000001010000", -- Line 1   Column 4017   Coefficient 72.07812500
   "010010000001010010", -- Line 1   Column 4018   Coefficient 72.08007813
   "010010000001010100", -- Line 1   Column 4019   Coefficient 72.08203125
   "010010000001010111", -- Line 1   Column 4020   Coefficient 72.08496094
   "010010000001011001", -- Line 1   Column 4021   Coefficient 72.08691406
   "010010000001011011", -- Line 1   Column 4022   Coefficient 72.08886719
   "010010000001011101", -- Line 1   Column 4023   Coefficient 72.09082031
   "010010000001011111", -- Line 1   Column 4024   Coefficient 72.09277344
   "010010000001100010", -- Line 1   Column 4025   Coefficient 72.09570313
   "010010000001100100", -- Line 1   Column 4026   Coefficient 72.09765625
   "010010000001100110", -- Line 1   Column 4027   Coefficient 72.09960938
   "010010000001101000", -- Line 1   Column 4028   Coefficient 72.10156250
   "010010000001101010", -- Line 1   Column 4029   Coefficient 72.10351563
   "010010000001101101", -- Line 1   Column 4030   Coefficient 72.10644531
   "010010000001101111", -- Line 1   Column 4031   Coefficient 72.10839844
   "010010000001110001", -- Line 1   Column 4032   Coefficient 72.11035156
   "010010000001110011", -- Line 1   Column 4033   Coefficient 72.11230469
   "010010000001110101", -- Line 1   Column 4034   Coefficient 72.11425781
   "010010000001111000", -- Line 1   Column 4035   Coefficient 72.11718750
   "010010000001111010", -- Line 1   Column 4036   Coefficient 72.11914063
   "010010000001111100", -- Line 1   Column 4037   Coefficient 72.12109375
   "010010000001111110", -- Line 1   Column 4038   Coefficient 72.12304688
   "010010000010000000", -- Line 1   Column 4039   Coefficient 72.12500000
   "010010000010000011", -- Line 1   Column 4040   Coefficient 72.12792969
   "010010000010000101", -- Line 1   Column 4041   Coefficient 72.12988281
   "010010000010000111", -- Line 1   Column 4042   Coefficient 72.13183594
   "010010000010001001", -- Line 1   Column 4043   Coefficient 72.13378906
   "010010000010001011", -- Line 1   Column 4044   Coefficient 72.13574219
   "010010000010001110", -- Line 1   Column 4045   Coefficient 72.13867188
   "010010000010010000", -- Line 1   Column 4046   Coefficient 72.14062500
   "010010000010010010", -- Line 1   Column 4047   Coefficient 72.14257813
   "010010000010010100", -- Line 1   Column 4048   Coefficient 72.14453125
   "010010000010010110", -- Line 1   Column 4049   Coefficient 72.14648438
   "010010000010011001", -- Line 1   Column 4050   Coefficient 72.14941406
   "010010000010011011", -- Line 1   Column 4051   Coefficient 72.15136719
   "010010000010011101", -- Line 1   Column 4052   Coefficient 72.15332031
   "010010000010011111", -- Line 1   Column 4053   Coefficient 72.15527344
   "010010000010100001", -- Line 1   Column 4054   Coefficient 72.15722656
   "010010000010100100", -- Line 1   Column 4055   Coefficient 72.16015625
   "010010000010100110", -- Line 1   Column 4056   Coefficient 72.16210938
   "010010000010101000", -- Line 1   Column 4057   Coefficient 72.16406250
   "010010000010101010", -- Line 1   Column 4058   Coefficient 72.16601563
   "010010000010101100", -- Line 1   Column 4059   Coefficient 72.16796875
   "010010000010101111", -- Line 1   Column 4060   Coefficient 72.17089844
   "010010000010110001", -- Line 1   Column 4061   Coefficient 72.17285156
   "010010000010110011", -- Line 1   Column 4062   Coefficient 72.17480469
   "010010000010110101", -- Line 1   Column 4063   Coefficient 72.17675781
   "010010000010110111", -- Line 1   Column 4064   Coefficient 72.17871094
   "010010000010111010", -- Line 1   Column 4065   Coefficient 72.18164063
   "010010000010111100", -- Line 1   Column 4066   Coefficient 72.18359375
   "010010000010111110", -- Line 1   Column 4067   Coefficient 72.18554688
   "010010000011000000", -- Line 1   Column 4068   Coefficient 72.18750000
   "010010000011000010", -- Line 1   Column 4069   Coefficient 72.18945313
   "010010000011000100", -- Line 1   Column 4070   Coefficient 72.19140625
   "010010000011000111", -- Line 1   Column 4071   Coefficient 72.19433594
   "010010000011001001", -- Line 1   Column 4072   Coefficient 72.19628906
   "010010000011001011", -- Line 1   Column 4073   Coefficient 72.19824219
   "010010000011001101", -- Line 1   Column 4074   Coefficient 72.20019531
   "010010000011001111", -- Line 1   Column 4075   Coefficient 72.20214844
   "010010000011010010", -- Line 1   Column 4076   Coefficient 72.20507813
   "010010000011010100", -- Line 1   Column 4077   Coefficient 72.20703125
   "010010000011010110", -- Line 1   Column 4078   Coefficient 72.20898438
   "010010000011011000", -- Line 1   Column 4079   Coefficient 72.21093750
   "010010000011011010", -- Line 1   Column 4080   Coefficient 72.21289063
   "010010000011011100", -- Line 1   Column 4081   Coefficient 72.21484375
   "010010000011011111", -- Line 1   Column 4082   Coefficient 72.21777344
   "010010000011100001", -- Line 1   Column 4083   Coefficient 72.21972656
   "010010000011100011", -- Line 1   Column 4084   Coefficient 72.22167969
   "010010000011100101", -- Line 1   Column 4085   Coefficient 72.22363281
   "010010000011100111", -- Line 1   Column 4086   Coefficient 72.22558594
   "010010000011101010", -- Line 1   Column 4087   Coefficient 72.22851563
   "010010000011101100", -- Line 1   Column 4088   Coefficient 72.23046875
   "010010000011101110", -- Line 1   Column 4089   Coefficient 72.23242188
   "010010000011110000", -- Line 1   Column 4090   Coefficient 72.23437500
   "010010000011110010", -- Line 1   Column 4091   Coefficient 72.23632813
   "010010000011110100", -- Line 1   Column 4092   Coefficient 72.23828125
   "010010000011110111", -- Line 1   Column 4093   Coefficient 72.24121094
   "010010000011111001", -- Line 1   Column 4094   Coefficient 72.24316406
   "010010000011111011", -- Line 1   Column 4095   Coefficient 72.24511719
   "010010000011111101" -- Line 1   Column 4096   Coefficient 72.24707031
);
begin
	process(clk)
	begin
	if(rising_edge(CLK)) then
		A <= rom(to_integer(unsigned(I)));
	end if;
	end process;
end ROM;
