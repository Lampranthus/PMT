-- DWT matrix coefficients
--
-- FI - UAQ
--
-- Electronica Avanzada III
--
-- Rene Romero Troncoso
--

library IEEE;
use IEEE.std_logic_1164.all;

entity ROM_DWT is
   port(
      I : in  std_logic_vector(11 downto 0);
      A : out std_logic_vector(17 downto 0)
      );
   end ROM_DWT;

architecture LUTable of ROM_DWT is
begin
   process(I)
   begin
      case I is
         -- Coefficient format 0.18
         when "000000000000" => A <= "000000000000001001"; -- Line 1   Column 1   Coefficient 0.00003433
         when "000000000001" => A <= "000000000000000011"; -- Line 1   Column 2   Coefficient 0.00001144
         when "000000000010" => A <= "111111111111001011"; -- Line 1   Column 3   Coefficient -0.00020218
         when "000000000011" => A <= "111111111110100110"; -- Line 1   Column 4   Coefficient -0.00034332
         when "000000000100" => A <= "111111111110010010"; -- Line 1   Column 5   Coefficient -0.00041962
         when "000000000101" => A <= "111111111111010011"; -- Line 1   Column 6   Coefficient -0.00017166
         when "000000000110" => A <= "000000000011111000"; -- Line 1   Column 7   Coefficient 0.00094604
         when "000000000111" => A <= "000000001000010011"; -- Line 1   Column 8   Coefficient 0.00202560
         when "000000001000" => A <= "000000001010110110"; -- Line 1   Column 9   Coefficient 0.00264740
         when "000000001001" => A <= "000000001101001100"; -- Line 1   Column 10   Coefficient 0.00321960
         when "000000001010" => A <= "000000001111111100"; -- Line 1   Column 11   Coefficient 0.00389099
         when "000000001011" => A <= "000000010000011000"; -- Line 1   Column 12   Coefficient 0.00399780
         when "000000001100" => A <= "000000001111000010"; -- Line 1   Column 13   Coefficient 0.00366974
         when "000000001101" => A <= "000000000111011010"; -- Line 1   Column 14   Coefficient 0.00180817
         when "000000001110" => A <= "111111110001010101"; -- Line 1   Column 15   Coefficient -0.00358200
         when "000000001111" => A <= "111111011001111001"; -- Line 1   Column 16   Coefficient -0.00930405
         when "000000010000" => A <= "111111000100111001"; -- Line 1   Column 17   Coefficient -0.01443100
         when "000000010001" => A <= "111110110001100001"; -- Line 1   Column 18   Coefficient -0.01916122
         when "000000010010" => A <= "111110100110010011"; -- Line 1   Column 19   Coefficient -0.02190018
         when "000000010011" => A <= "111110011011111010"; -- Line 1   Column 20   Coefficient -0.02443695
         when "000000010100" => A <= "111110010000110000"; -- Line 1   Column 21   Coefficient -0.02716064
         when "000000010101" => A <= "111110000101010011"; -- Line 1   Column 22   Coefficient -0.02995682
         when "000000010110" => A <= "111101110100001010"; -- Line 1   Column 23   Coefficient -0.03414154
         when "000000010111" => A <= "111101100110110000"; -- Line 1   Column 24   Coefficient -0.03741455
         when "000000011000" => A <= "111101100010101111"; -- Line 1   Column 25   Coefficient -0.03839493
         when "000000011001" => A <= "111101100010001110"; -- Line 1   Column 26   Coefficient -0.03852081
         when "000000011010" => A <= "111101100000101101"; -- Line 1   Column 27   Coefficient -0.03889084
         when "000000011011" => A <= "111101101011101110"; -- Line 1   Column 28   Coefficient -0.03620148
         when "000000011100" => A <= "111110000010011110"; -- Line 1   Column 29   Coefficient -0.03064728
         when "000000011101" => A <= "111110110101100100"; -- Line 1   Column 30   Coefficient -0.01817322
         when "000000011110" => A <= "000000100101011001"; -- Line 1   Column 31   Coefficient 0.00912857
         when "000000011111" => A <= "000010011110111100"; -- Line 1   Column 32   Coefficient 0.03880310
         when "000000100000" => A <= "000100010010000101"; -- Line 1   Column 33   Coefficient 0.06691360
         when "000000100001" => A <= "000110000101110011"; -- Line 1   Column 34   Coefficient 0.09516525
         when "000000100010" => A <= "000111100110110001"; -- Line 1   Column 35   Coefficient 0.11883926
         when "000000100011" => A <= "001001000110101001"; -- Line 1   Column 36   Coefficient 0.14224625
         when "000000100100" => A <= "001010101100000111"; -- Line 1   Column 37   Coefficient 0.16701889
         when "000000100101" => A <= "001100001011101000"; -- Line 1   Column 38   Coefficient 0.19033813
         when "000000100110" => A <= "001101100011111111"; -- Line 1   Column 39   Coefficient 0.21191025
         when "000000100111" => A <= "001110110101010100"; -- Line 1   Column 40   Coefficient 0.23176575
         when "000000101000" => A <= "001111111010100001"; -- Line 1   Column 41   Coefficient 0.24866104
         when "000000101001" => A <= "010000111010100101"; -- Line 1   Column 42   Coefficient 0.26430130
         when "000000101010" => A <= "010010000001100011"; -- Line 1   Column 43   Coefficient 0.28162766
         when "000000101011" => A <= "010010110100110100"; -- Line 1   Column 44   Coefficient 0.29414368
         when "000000101100" => A <= "010011010010100110"; -- Line 1   Column 45   Coefficient 0.30141449
         when "000000101101" => A <= "010011000101100111"; -- Line 1   Column 46   Coefficient 0.29824448
         when "000000101110" => A <= "010001011110001011"; -- Line 1   Column 47   Coefficient 0.27299118
         when "000000101111" => A <= "001111100101110011"; -- Line 1   Column 48   Coefficient 0.24360275
         when "000000110000" => A <= "001101110100101001"; -- Line 1   Column 49   Coefficient 0.21597672
         when "000000110001" => A <= "001011111101111010"; -- Line 1   Column 50   Coefficient 0.18698883
         when "000000110010" => A <= "001010011001111000"; -- Line 1   Column 51   Coefficient 0.16256714
         when "000000110011" => A <= "001000110101000000"; -- Line 1   Column 52   Coefficient 0.13793945
         when "000000110100" => A <= "000111000101010101"; -- Line 1   Column 53   Coefficient 0.11067581
         when "000000110101" => A <= "000101100000010101"; -- Line 1   Column 54   Coefficient 0.08601761
         when "000000110110" => A <= "000100010011001101"; -- Line 1   Column 55   Coefficient 0.06718826
         when "000000110111" => A <= "000011001010010011"; -- Line 1   Column 56   Coefficient 0.04938889
         when "000000111000" => A <= "000010000100001011"; -- Line 1   Column 57   Coefficient 0.03226852
         when "000000111001" => A <= "000000111110100110"; -- Line 1   Column 58   Coefficient 0.01528168
         when "000000111010" => A <= "111111101010001000"; -- Line 1   Column 59   Coefficient -0.00534058
         when "000000111011" => A <= "111110100000101100"; -- Line 1   Column 60   Coefficient -0.02326965
         when "000000111100" => A <= "111101100111001110"; -- Line 1   Column 61   Coefficient -0.03730011
         when "000000111101" => A <= "111101000110110001"; -- Line 1   Column 62   Coefficient -0.04522324
         when "000000111110" => A <= "111101011101101101"; -- Line 1   Column 63   Coefficient -0.03962326
         when "000000111111" => A <= "111101111110110001"; -- Line 1   Column 64   Coefficient -0.03155136
         when "000001000000" => A <= "111110011010010101"; -- Line 1   Column 65   Coefficient -0.02482224
         when "000001000001" => A <= "111110111010000001"; -- Line 1   Column 66   Coefficient -0.01708603
         when "000001000010" => A <= "111111010000101110"; -- Line 1   Column 67   Coefficient -0.01154327
         when "000001000011" => A <= "111111100111100010"; -- Line 1   Column 68   Coefficient -0.00597382
         when "000001000100" => A <= "000000000100100100"; -- Line 1   Column 69   Coefficient 0.00111389
         when "000001000101" => A <= "000000011000110111"; -- Line 1   Column 70   Coefficient 0.00606918
         when "000001000110" => A <= "000000010111101010"; -- Line 1   Column 71   Coefficient 0.00577545
         when "000001000111" => A <= "000000010100111001"; -- Line 1   Column 72   Coefficient 0.00510025
         when "000001001000" => A <= "000000010100110111"; -- Line 1   Column 73   Coefficient 0.00509262
         when "000001001001" => A <= "000000010110010000"; -- Line 1   Column 74   Coefficient 0.00543213
         when "000001001010" => A <= "000000100010100100"; -- Line 1   Column 75   Coefficient 0.00843811
         when "000001001011" => A <= "000000101101010111"; -- Line 1   Column 76   Coefficient 0.01107407
         when "000001001100" => A <= "000000110010101110"; -- Line 1   Column 77   Coefficient 0.01238251
         when "000001001101" => A <= "000000110100010110"; -- Line 1   Column 78   Coefficient 0.01277924
         when "000001001110" => A <= "000000101011110101"; -- Line 1   Column 79   Coefficient 0.01070023
         when "000001001111" => A <= "000000100001110011"; -- Line 1   Column 80   Coefficient 0.00825119
         when "000001010000" => A <= "000000011001110100"; -- Line 1   Column 81   Coefficient 0.00630188
         when "000001010001" => A <= "000000010001001000"; -- Line 1   Column 82   Coefficient 0.00418091
         when "000001010010" => A <= "000000001001011000"; -- Line 1   Column 83   Coefficient 0.00228882
         when "000001010011" => A <= "000000000010010011"; -- Line 1   Column 84   Coefficient 0.00056076
         when "000001010100" => A <= "111111111010111001"; -- Line 1   Column 85   Coefficient -0.00124741
         when "000001010101" => A <= "111111110110011111"; -- Line 1   Column 86   Coefficient -0.00232315
         when "000001010110" => A <= "111111111001000110"; -- Line 1   Column 87   Coefficient -0.00168610
         when "000001010111" => A <= "111111111100011110"; -- Line 1   Column 88   Coefficient -0.00086212
         when "000001011000" => A <= "111111111110110111"; -- Line 1   Column 89   Coefficient -0.00027847
         when "000001011001" => A <= "000000000001001011"; -- Line 1   Column 90   Coefficient 0.00028610
         when "000001011010" => A <= "000000000001001000"; -- Line 1   Column 91   Coefficient 0.00027466
         when "000001011011" => A <= "000000000001000010"; -- Line 1   Column 92   Coefficient 0.00025177
         when "000001011100" => A <= "000000000001111110"; -- Line 1   Column 93   Coefficient 0.00048065
         when "000001011101" => A <= "000000000010010101"; -- Line 1   Column 94   Coefficient 0.00056839
         when "000001011110" => A <= "000000000001100101"; -- Line 1   Column 95   Coefficient 0.00038528
         when "000001011111" => A <= "000000000000110011"; -- Line 1   Column 96   Coefficient 0.00019455
         when "000001100000" => A <= "000000000000000111"; -- Line 1   Column 97   Coefficient 0.00002670
         when "000001100001" => A <= "111111111111100110"; -- Line 1   Column 98   Coefficient -0.00009918
         when "000001100010" => A <= "111111111111110100"; -- Line 1   Column 99   Coefficient -0.00004578
         when "000001100011" => A <= "000000000000000011"; -- Line 1   Column 100   Coefficient 0.00001144
         when "000001100100" => A <= "000000000000000100"; -- Line 1   Column 101   Coefficient 0.00001526
         when "000001100101" => A <= "000000000000000110"; -- Line 1   Column 102   Coefficient 0.00002289
         when "000001100110" => A <= "000000000000000011"; -- Line 1   Column 103   Coefficient 0.00001144
         when "000001100111" => A <= "111111111111111111"; -- Line 1   Column 104   Coefficient -0.00000381
         when "000001101000" => A <= "000000000000000000"; -- Line 1   Column 105   Coefficient 0.00000000
         when "000001101001" => A <= "000000000000000000"; -- Line 1   Column 106   Coefficient 0.00000000
         when "000001101010" => A <= "000000000000000000"; -- Line 1   Column 107   Coefficient 0.00000000
         when "000001101011" => A <= "000000000000000000"; -- Line 1   Column 108   Coefficient 0.00000000
         when "000001101100" => A <= "000000000000000000"; -- Line 1   Column 109   Coefficient 0.00000000
         when "000001101101" => A <= "000000000000000000"; -- Line 1   Column 110   Coefficient 0.00000000
         when "000001101110" => A <= "000000000000000000"; -- Line 1   Column 111   Coefficient 0.00000000
         when "000001101111" => A <= "000000000000000000"; -- Line 1   Column 112   Coefficient 0.00000000
         when "000001110000" => A <= "000000000000000000"; -- Line 1   Column 113   Coefficient 0.00000000
         when "000001110001" => A <= "000000000000000000"; -- Line 1   Column 114   Coefficient 0.00000000
         when "000001110010" => A <= "000000000000000000"; -- Line 1   Column 115   Coefficient 0.00000000
         when "000001110011" => A <= "000000000000000000"; -- Line 1   Column 116   Coefficient 0.00000000
         when "000001110100" => A <= "000000000000000000"; -- Line 1   Column 117   Coefficient 0.00000000
         when "000001110101" => A <= "000000000000000000"; -- Line 1   Column 118   Coefficient 0.00000000
         when "000001110110" => A <= "000000000000000000"; -- Line 1   Column 119   Coefficient 0.00000000
         when "000001110111" => A <= "000000000000000000"; -- Line 1   Column 120   Coefficient 0.00000000
         when "000001111000" => A <= "000000000000000000"; -- Line 1   Column 121   Coefficient 0.00000000
         when "000001111001" => A <= "000000000000000000"; -- Line 1   Column 122   Coefficient 0.00000000
         when "000001111010" => A <= "000000000000000000"; -- Line 1   Column 123   Coefficient 0.00000000
         when "000001111011" => A <= "000000000000000000"; -- Line 1   Column 124   Coefficient 0.00000000
         when "000001111100" => A <= "000000000000000000"; -- Line 1   Column 125   Coefficient 0.00000000
         when "000001111101" => A <= "000000000000000000"; -- Line 1   Column 126   Coefficient 0.00000000
         when "000001111110" => A <= "000000000000000000"; -- Line 1   Column 127   Coefficient 0.00000000
         when "000001111111" => A <= "000000000000000000"; -- Line 1   Column 128   Coefficient 0.00000000
         when "000010000000" => A <= "000000000000000000"; -- Line 1   Column 129   Coefficient 0.00000000
         when "000010000001" => A <= "000000000000000000"; -- Line 1   Column 130   Coefficient 0.00000000
         when "000010000010" => A <= "000000000000000000"; -- Line 1   Column 131   Coefficient 0.00000000
         when "000010000011" => A <= "000000000000000000"; -- Line 1   Column 132   Coefficient 0.00000000
         when "000010000100" => A <= "000000000000000000"; -- Line 1   Column 133   Coefficient 0.00000000
         when "000010000101" => A <= "000000000000000000"; -- Line 1   Column 134   Coefficient 0.00000000
         when "000010000110" => A <= "000000000000000000"; -- Line 1   Column 135   Coefficient 0.00000000
         when "000010000111" => A <= "000000000000000000"; -- Line 1   Column 136   Coefficient 0.00000000
         when "000010001000" => A <= "000000000000000000"; -- Line 1   Column 137   Coefficient 0.00000000
         when "000010001001" => A <= "000000000000000000"; -- Line 1   Column 138   Coefficient 0.00000000
         when "000010001010" => A <= "000000000000000000"; -- Line 1   Column 139   Coefficient 0.00000000
         when "000010001011" => A <= "000000000000000000"; -- Line 1   Column 140   Coefficient 0.00000000
         when "000010001100" => A <= "000000000000000000"; -- Line 1   Column 141   Coefficient 0.00000000
         when "000010001101" => A <= "000000000000000000"; -- Line 1   Column 142   Coefficient 0.00000000
         when "000010001110" => A <= "000000000000000000"; -- Line 1   Column 143   Coefficient 0.00000000
         when "000010001111" => A <= "000000000000000000"; -- Line 1   Column 144   Coefficient 0.00000000
         when "000010010000" => A <= "000000000000000000"; -- Line 1   Column 145   Coefficient 0.00000000
         when "000010010001" => A <= "000000000000000000"; -- Line 1   Column 146   Coefficient 0.00000000
         when "000010010010" => A <= "000000000000000000"; -- Line 1   Column 147   Coefficient 0.00000000
         when "000010010011" => A <= "000000000000000000"; -- Line 1   Column 148   Coefficient 0.00000000
         when "000010010100" => A <= "000000000000000000"; -- Line 1   Column 149   Coefficient 0.00000000
         when "000010010101" => A <= "000000000000000000"; -- Line 1   Column 150   Coefficient 0.00000000
         when "000010010110" => A <= "000000000000000000"; -- Line 1   Column 151   Coefficient 0.00000000
         when "000010010111" => A <= "000000000000000000"; -- Line 1   Column 152   Coefficient 0.00000000
         when "000010011000" => A <= "000000000000000000"; -- Line 1   Column 153   Coefficient 0.00000000
         when "000010011001" => A <= "000000000000000000"; -- Line 1   Column 154   Coefficient 0.00000000
         when "000010011010" => A <= "000000000000000000"; -- Line 1   Column 155   Coefficient 0.00000000
         when "000010011011" => A <= "000000000000000000"; -- Line 1   Column 156   Coefficient 0.00000000
         when "000010011100" => A <= "000000000000000000"; -- Line 1   Column 157   Coefficient 0.00000000
         when "000010011101" => A <= "000000000000000000"; -- Line 1   Column 158   Coefficient 0.00000000
         when "000010011110" => A <= "000000000000000000"; -- Line 1   Column 159   Coefficient 0.00000000
         when "000010011111" => A <= "000000000000000000"; -- Line 1   Column 160   Coefficient 0.00000000
         when "000010100000" => A <= "000000000000000000"; -- Line 1   Column 161   Coefficient 0.00000000
         when "000010100001" => A <= "000000000000000000"; -- Line 1   Column 162   Coefficient 0.00000000
         when "000010100010" => A <= "000000000000000000"; -- Line 1   Column 163   Coefficient 0.00000000
         when "000010100011" => A <= "000000000000000000"; -- Line 1   Column 164   Coefficient 0.00000000
         when "000010100100" => A <= "000000000000000000"; -- Line 1   Column 165   Coefficient 0.00000000
         when "000010100101" => A <= "000000000000000000"; -- Line 1   Column 166   Coefficient 0.00000000
         when "000010100110" => A <= "000000000000000000"; -- Line 1   Column 167   Coefficient 0.00000000
         when "000010100111" => A <= "000000000000000000"; -- Line 1   Column 168   Coefficient 0.00000000
         when "000010101000" => A <= "000000000000000000"; -- Line 1   Column 169   Coefficient 0.00000000
         when "000010101001" => A <= "000000000000000000"; -- Line 1   Column 170   Coefficient 0.00000000
         when "000010101010" => A <= "000000000000000000"; -- Line 1   Column 171   Coefficient 0.00000000
         when "000010101011" => A <= "000000000000000000"; -- Line 1   Column 172   Coefficient 0.00000000
         when "000010101100" => A <= "000000000000000000"; -- Line 1   Column 173   Coefficient 0.00000000
         when "000010101101" => A <= "000000000000000000"; -- Line 1   Column 174   Coefficient 0.00000000
         when "000010101110" => A <= "000000000000000000"; -- Line 1   Column 175   Coefficient 0.00000000
         when "000010101111" => A <= "000000000000000000"; -- Line 1   Column 176   Coefficient 0.00000000
         when "000010110000" => A <= "000000000000000000"; -- Line 1   Column 177   Coefficient 0.00000000
         when "000010110001" => A <= "000000000000000000"; -- Line 1   Column 178   Coefficient 0.00000000
         when "000010110010" => A <= "000000000000000000"; -- Line 1   Column 179   Coefficient 0.00000000
         when "000010110011" => A <= "000000000000000000"; -- Line 1   Column 180   Coefficient 0.00000000
         when "000010110100" => A <= "000000000000000000"; -- Line 1   Column 181   Coefficient 0.00000000
         when "000010110101" => A <= "000000000000000000"; -- Line 1   Column 182   Coefficient 0.00000000
         when "000010110110" => A <= "000000000000000000"; -- Line 1   Column 183   Coefficient 0.00000000
         when "000010110111" => A <= "000000000000000000"; -- Line 1   Column 184   Coefficient 0.00000000
         when "000010111000" => A <= "000000000000000000"; -- Line 1   Column 185   Coefficient 0.00000000
         when "000010111001" => A <= "000000000000000000"; -- Line 1   Column 186   Coefficient 0.00000000
         when "000010111010" => A <= "000000000000000000"; -- Line 1   Column 187   Coefficient 0.00000000
         when "000010111011" => A <= "000000000000000000"; -- Line 1   Column 188   Coefficient 0.00000000
         when "000010111100" => A <= "000000000000000000"; -- Line 1   Column 189   Coefficient 0.00000000
         when "000010111101" => A <= "000000000000000000"; -- Line 1   Column 190   Coefficient 0.00000000
         when "000010111110" => A <= "000000000000000000"; -- Line 1   Column 191   Coefficient 0.00000000
         when "000010111111" => A <= "000000000000000000"; -- Line 1   Column 192   Coefficient 0.00000000
         when "000011000000" => A <= "000000000000000000"; -- Line 1   Column 193   Coefficient 0.00000000
         when "000011000001" => A <= "000000000000000000"; -- Line 1   Column 194   Coefficient 0.00000000
         when "000011000010" => A <= "000000000000000000"; -- Line 1   Column 195   Coefficient 0.00000000
         when "000011000011" => A <= "000000000000000000"; -- Line 1   Column 196   Coefficient 0.00000000
         when "000011000100" => A <= "000000000000000000"; -- Line 1   Column 197   Coefficient 0.00000000
         when "000011000101" => A <= "000000000000000000"; -- Line 1   Column 198   Coefficient 0.00000000
         when "000011000110" => A <= "000000000000000000"; -- Line 1   Column 199   Coefficient 0.00000000
         when "000011000111" => A <= "000000000000000000"; -- Line 1   Column 200   Coefficient 0.00000000
         when "000011001000" => A <= "000000000000000000"; -- Line 1   Column 201   Coefficient 0.00000000
         when "000011001001" => A <= "000000000000000000"; -- Line 1   Column 202   Coefficient 0.00000000
         when "000011001010" => A <= "000000000000000000"; -- Line 1   Column 203   Coefficient 0.00000000
         when "000011001011" => A <= "000000000000000000"; -- Line 1   Column 204   Coefficient 0.00000000
         when "000011001100" => A <= "000000000000000000"; -- Line 1   Column 205   Coefficient 0.00000000
         when "000011001101" => A <= "000000000000000000"; -- Line 1   Column 206   Coefficient 0.00000000
         when "000011001110" => A <= "000000000000000000"; -- Line 1   Column 207   Coefficient 0.00000000
         when "000011001111" => A <= "000000000000000000"; -- Line 1   Column 208   Coefficient 0.00000000
         when "000011010000" => A <= "000000000000000000"; -- Line 1   Column 209   Coefficient 0.00000000
         when "000011010001" => A <= "000000000000000000"; -- Line 1   Column 210   Coefficient 0.00000000
         when "000011010010" => A <= "000000000000000000"; -- Line 1   Column 211   Coefficient 0.00000000
         when "000011010011" => A <= "000000000000000000"; -- Line 1   Column 212   Coefficient 0.00000000
         when "000011010100" => A <= "000000000000000000"; -- Line 1   Column 213   Coefficient 0.00000000
         when "000011010101" => A <= "000000000000000000"; -- Line 1   Column 214   Coefficient 0.00000000
         when "000011010110" => A <= "000000000000000000"; -- Line 1   Column 215   Coefficient 0.00000000
         when "000011010111" => A <= "000000000000000000"; -- Line 1   Column 216   Coefficient 0.00000000
         when "000011011000" => A <= "000000000000000000"; -- Line 1   Column 217   Coefficient 0.00000000
         when "000011011001" => A <= "000000000000000000"; -- Line 1   Column 218   Coefficient 0.00000000
         when "000011011010" => A <= "000000000000000000"; -- Line 1   Column 219   Coefficient 0.00000000
         when "000011011011" => A <= "000000000000000000"; -- Line 1   Column 220   Coefficient 0.00000000
         when "000011011100" => A <= "000000000000000000"; -- Line 1   Column 221   Coefficient 0.00000000
         when "000011011101" => A <= "000000000000000000"; -- Line 1   Column 222   Coefficient 0.00000000
         when "000011011110" => A <= "000000000000000000"; -- Line 1   Column 223   Coefficient 0.00000000
         when "000011011111" => A <= "000000000000000000"; -- Line 1   Column 224   Coefficient 0.00000000
         when "000011100000" => A <= "000000000000000000"; -- Line 1   Column 225   Coefficient 0.00000000
         when "000011100001" => A <= "000000000000000000"; -- Line 1   Column 226   Coefficient 0.00000000
         when "000011100010" => A <= "000000000000000000"; -- Line 1   Column 227   Coefficient 0.00000000
         when "000011100011" => A <= "000000000000000000"; -- Line 1   Column 228   Coefficient 0.00000000
         when "000011100100" => A <= "000000000000000000"; -- Line 1   Column 229   Coefficient 0.00000000
         when "000011100101" => A <= "000000000000000000"; -- Line 1   Column 230   Coefficient 0.00000000
         when "000011100110" => A <= "000000000000000000"; -- Line 1   Column 231   Coefficient 0.00000000
         when "000011100111" => A <= "000000000000000000"; -- Line 1   Column 232   Coefficient 0.00000000
         when "000011101000" => A <= "000000000000000000"; -- Line 1   Column 233   Coefficient 0.00000000
         when "000011101001" => A <= "000000000000000000"; -- Line 1   Column 234   Coefficient 0.00000000
         when "000011101010" => A <= "000000000000000000"; -- Line 1   Column 235   Coefficient 0.00000000
         when "000011101011" => A <= "000000000000000000"; -- Line 1   Column 236   Coefficient 0.00000000
         when "000011101100" => A <= "000000000000000000"; -- Line 1   Column 237   Coefficient 0.00000000
         when "000011101101" => A <= "000000000000000000"; -- Line 1   Column 238   Coefficient 0.00000000
         when "000011101110" => A <= "000000000000000000"; -- Line 1   Column 239   Coefficient 0.00000000
         when "000011101111" => A <= "000000000000000000"; -- Line 1   Column 240   Coefficient 0.00000000
         when "000011110000" => A <= "000000000000000000"; -- Line 1   Column 241   Coefficient 0.00000000
         when "000011110001" => A <= "000000000000000000"; -- Line 1   Column 242   Coefficient 0.00000000
         when "000011110010" => A <= "000000000000000000"; -- Line 1   Column 243   Coefficient 0.00000000
         when "000011110011" => A <= "000000000000000000"; -- Line 1   Column 244   Coefficient 0.00000000
         when "000011110100" => A <= "000000000000000000"; -- Line 1   Column 245   Coefficient 0.00000000
         when "000011110101" => A <= "000000000000000000"; -- Line 1   Column 246   Coefficient 0.00000000
         when "000011110110" => A <= "000000000000000000"; -- Line 1   Column 247   Coefficient 0.00000000
         when "000011110111" => A <= "000000000000000000"; -- Line 1   Column 248   Coefficient 0.00000000
         when "000011111000" => A <= "000000000000000000"; -- Line 1   Column 249   Coefficient 0.00000000
         when "000011111001" => A <= "000000000000000000"; -- Line 1   Column 250   Coefficient 0.00000000
         when "000011111010" => A <= "000000000000000000"; -- Line 1   Column 251   Coefficient 0.00000000
         when "000011111011" => A <= "000000000000000000"; -- Line 1   Column 252   Coefficient 0.00000000
         when "000011111100" => A <= "000000000000000000"; -- Line 1   Column 253   Coefficient 0.00000000
         when "000011111101" => A <= "000000000000000000"; -- Line 1   Column 254   Coefficient 0.00000000
         when "000011111110" => A <= "000000000000000000"; -- Line 1   Column 255   Coefficient 0.00000000
         when "000011111111" => A <= "000000000000000000"; -- Line 1   Column 256   Coefficient 0.00000000
         when "000100000000" => A <= "000000000000000000"; -- Line 2   Column 1   Coefficient 0.00000000
         when "000100000001" => A <= "000000000000000000"; -- Line 2   Column 2   Coefficient 0.00000000
         when "000100000010" => A <= "000000000000000000"; -- Line 2   Column 3   Coefficient 0.00000000
         when "000100000011" => A <= "000000000000000000"; -- Line 2   Column 4   Coefficient 0.00000000
         when "000100000100" => A <= "000000000000000000"; -- Line 2   Column 5   Coefficient 0.00000000
         when "000100000101" => A <= "000000000000000000"; -- Line 2   Column 6   Coefficient 0.00000000
         when "000100000110" => A <= "000000000000000000"; -- Line 2   Column 7   Coefficient 0.00000000
         when "000100000111" => A <= "000000000000000000"; -- Line 2   Column 8   Coefficient 0.00000000
         when "000100001000" => A <= "000000000000000000"; -- Line 2   Column 9   Coefficient 0.00000000
         when "000100001001" => A <= "000000000000000000"; -- Line 2   Column 10   Coefficient 0.00000000
         when "000100001010" => A <= "000000000000000000"; -- Line 2   Column 11   Coefficient 0.00000000
         when "000100001011" => A <= "000000000000000000"; -- Line 2   Column 12   Coefficient 0.00000000
         when "000100001100" => A <= "000000000000000000"; -- Line 2   Column 13   Coefficient 0.00000000
         when "000100001101" => A <= "000000000000000000"; -- Line 2   Column 14   Coefficient 0.00000000
         when "000100001110" => A <= "000000000000000000"; -- Line 2   Column 15   Coefficient 0.00000000
         when "000100001111" => A <= "000000000000000000"; -- Line 2   Column 16   Coefficient 0.00000000
         when "000100010000" => A <= "000000000000001001"; -- Line 2   Column 17   Coefficient 0.00003433
         when "000100010001" => A <= "000000000000000011"; -- Line 2   Column 18   Coefficient 0.00001144
         when "000100010010" => A <= "111111111111001011"; -- Line 2   Column 19   Coefficient -0.00020218
         when "000100010011" => A <= "111111111110100110"; -- Line 2   Column 20   Coefficient -0.00034332
         when "000100010100" => A <= "111111111110010010"; -- Line 2   Column 21   Coefficient -0.00041962
         when "000100010101" => A <= "111111111111010011"; -- Line 2   Column 22   Coefficient -0.00017166
         when "000100010110" => A <= "000000000011111000"; -- Line 2   Column 23   Coefficient 0.00094604
         when "000100010111" => A <= "000000001000010011"; -- Line 2   Column 24   Coefficient 0.00202560
         when "000100011000" => A <= "000000001010110110"; -- Line 2   Column 25   Coefficient 0.00264740
         when "000100011001" => A <= "000000001101001100"; -- Line 2   Column 26   Coefficient 0.00321960
         when "000100011010" => A <= "000000001111111100"; -- Line 2   Column 27   Coefficient 0.00389099
         when "000100011011" => A <= "000000010000011000"; -- Line 2   Column 28   Coefficient 0.00399780
         when "000100011100" => A <= "000000001111000010"; -- Line 2   Column 29   Coefficient 0.00366974
         when "000100011101" => A <= "000000000111011010"; -- Line 2   Column 30   Coefficient 0.00180817
         when "000100011110" => A <= "111111110001010101"; -- Line 2   Column 31   Coefficient -0.00358200
         when "000100011111" => A <= "111111011001111001"; -- Line 2   Column 32   Coefficient -0.00930405
         when "000100100000" => A <= "111111000100111001"; -- Line 2   Column 33   Coefficient -0.01443100
         when "000100100001" => A <= "111110110001100001"; -- Line 2   Column 34   Coefficient -0.01916122
         when "000100100010" => A <= "111110100110010011"; -- Line 2   Column 35   Coefficient -0.02190018
         when "000100100011" => A <= "111110011011111010"; -- Line 2   Column 36   Coefficient -0.02443695
         when "000100100100" => A <= "111110010000110000"; -- Line 2   Column 37   Coefficient -0.02716064
         when "000100100101" => A <= "111110000101010011"; -- Line 2   Column 38   Coefficient -0.02995682
         when "000100100110" => A <= "111101110100001010"; -- Line 2   Column 39   Coefficient -0.03414154
         when "000100100111" => A <= "111101100110110000"; -- Line 2   Column 40   Coefficient -0.03741455
         when "000100101000" => A <= "111101100010101111"; -- Line 2   Column 41   Coefficient -0.03839493
         when "000100101001" => A <= "111101100010001110"; -- Line 2   Column 42   Coefficient -0.03852081
         when "000100101010" => A <= "111101100000101101"; -- Line 2   Column 43   Coefficient -0.03889084
         when "000100101011" => A <= "111101101011101110"; -- Line 2   Column 44   Coefficient -0.03620148
         when "000100101100" => A <= "111110000010011110"; -- Line 2   Column 45   Coefficient -0.03064728
         when "000100101101" => A <= "111110110101100100"; -- Line 2   Column 46   Coefficient -0.01817322
         when "000100101110" => A <= "000000100101011001"; -- Line 2   Column 47   Coefficient 0.00912857
         when "000100101111" => A <= "000010011110111100"; -- Line 2   Column 48   Coefficient 0.03880310
         when "000100110000" => A <= "000100010010000101"; -- Line 2   Column 49   Coefficient 0.06691360
         when "000100110001" => A <= "000110000101110011"; -- Line 2   Column 50   Coefficient 0.09516525
         when "000100110010" => A <= "000111100110110001"; -- Line 2   Column 51   Coefficient 0.11883926
         when "000100110011" => A <= "001001000110101001"; -- Line 2   Column 52   Coefficient 0.14224625
         when "000100110100" => A <= "001010101100000111"; -- Line 2   Column 53   Coefficient 0.16701889
         when "000100110101" => A <= "001100001011101000"; -- Line 2   Column 54   Coefficient 0.19033813
         when "000100110110" => A <= "001101100011111111"; -- Line 2   Column 55   Coefficient 0.21191025
         when "000100110111" => A <= "001110110101010100"; -- Line 2   Column 56   Coefficient 0.23176575
         when "000100111000" => A <= "001111111010100001"; -- Line 2   Column 57   Coefficient 0.24866104
         when "000100111001" => A <= "010000111010100101"; -- Line 2   Column 58   Coefficient 0.26430130
         when "000100111010" => A <= "010010000001100011"; -- Line 2   Column 59   Coefficient 0.28162766
         when "000100111011" => A <= "010010110100110100"; -- Line 2   Column 60   Coefficient 0.29414368
         when "000100111100" => A <= "010011010010100110"; -- Line 2   Column 61   Coefficient 0.30141449
         when "000100111101" => A <= "010011000101100111"; -- Line 2   Column 62   Coefficient 0.29824448
         when "000100111110" => A <= "010001011110001011"; -- Line 2   Column 63   Coefficient 0.27299118
         when "000100111111" => A <= "001111100101110011"; -- Line 2   Column 64   Coefficient 0.24360275
         when "000101000000" => A <= "001101110100101001"; -- Line 2   Column 65   Coefficient 0.21597672
         when "000101000001" => A <= "001011111101111010"; -- Line 2   Column 66   Coefficient 0.18698883
         when "000101000010" => A <= "001010011001111000"; -- Line 2   Column 67   Coefficient 0.16256714
         when "000101000011" => A <= "001000110101000000"; -- Line 2   Column 68   Coefficient 0.13793945
         when "000101000100" => A <= "000111000101010101"; -- Line 2   Column 69   Coefficient 0.11067581
         when "000101000101" => A <= "000101100000010101"; -- Line 2   Column 70   Coefficient 0.08601761
         when "000101000110" => A <= "000100010011001101"; -- Line 2   Column 71   Coefficient 0.06718826
         when "000101000111" => A <= "000011001010010011"; -- Line 2   Column 72   Coefficient 0.04938889
         when "000101001000" => A <= "000010000100001011"; -- Line 2   Column 73   Coefficient 0.03226852
         when "000101001001" => A <= "000000111110100110"; -- Line 2   Column 74   Coefficient 0.01528168
         when "000101001010" => A <= "111111101010001000"; -- Line 2   Column 75   Coefficient -0.00534058
         when "000101001011" => A <= "111110100000101100"; -- Line 2   Column 76   Coefficient -0.02326965
         when "000101001100" => A <= "111101100111001110"; -- Line 2   Column 77   Coefficient -0.03730011
         when "000101001101" => A <= "111101000110110001"; -- Line 2   Column 78   Coefficient -0.04522324
         when "000101001110" => A <= "111101011101101101"; -- Line 2   Column 79   Coefficient -0.03962326
         when "000101001111" => A <= "111101111110110001"; -- Line 2   Column 80   Coefficient -0.03155136
         when "000101010000" => A <= "111110011010010101"; -- Line 2   Column 81   Coefficient -0.02482224
         when "000101010001" => A <= "111110111010000001"; -- Line 2   Column 82   Coefficient -0.01708603
         when "000101010010" => A <= "111111010000101110"; -- Line 2   Column 83   Coefficient -0.01154327
         when "000101010011" => A <= "111111100111100010"; -- Line 2   Column 84   Coefficient -0.00597382
         when "000101010100" => A <= "000000000100100100"; -- Line 2   Column 85   Coefficient 0.00111389
         when "000101010101" => A <= "000000011000110111"; -- Line 2   Column 86   Coefficient 0.00606918
         when "000101010110" => A <= "000000010111101010"; -- Line 2   Column 87   Coefficient 0.00577545
         when "000101010111" => A <= "000000010100111001"; -- Line 2   Column 88   Coefficient 0.00510025
         when "000101011000" => A <= "000000010100110111"; -- Line 2   Column 89   Coefficient 0.00509262
         when "000101011001" => A <= "000000010110010000"; -- Line 2   Column 90   Coefficient 0.00543213
         when "000101011010" => A <= "000000100010100100"; -- Line 2   Column 91   Coefficient 0.00843811
         when "000101011011" => A <= "000000101101010111"; -- Line 2   Column 92   Coefficient 0.01107407
         when "000101011100" => A <= "000000110010101110"; -- Line 2   Column 93   Coefficient 0.01238251
         when "000101011101" => A <= "000000110100010110"; -- Line 2   Column 94   Coefficient 0.01277924
         when "000101011110" => A <= "000000101011110101"; -- Line 2   Column 95   Coefficient 0.01070023
         when "000101011111" => A <= "000000100001110011"; -- Line 2   Column 96   Coefficient 0.00825119
         when "000101100000" => A <= "000000011001110100"; -- Line 2   Column 97   Coefficient 0.00630188
         when "000101100001" => A <= "000000010001001000"; -- Line 2   Column 98   Coefficient 0.00418091
         when "000101100010" => A <= "000000001001011000"; -- Line 2   Column 99   Coefficient 0.00228882
         when "000101100011" => A <= "000000000010010011"; -- Line 2   Column 100   Coefficient 0.00056076
         when "000101100100" => A <= "111111111010111001"; -- Line 2   Column 101   Coefficient -0.00124741
         when "000101100101" => A <= "111111110110011111"; -- Line 2   Column 102   Coefficient -0.00232315
         when "000101100110" => A <= "111111111001000110"; -- Line 2   Column 103   Coefficient -0.00168610
         when "000101100111" => A <= "111111111100011110"; -- Line 2   Column 104   Coefficient -0.00086212
         when "000101101000" => A <= "111111111110110111"; -- Line 2   Column 105   Coefficient -0.00027847
         when "000101101001" => A <= "000000000001001011"; -- Line 2   Column 106   Coefficient 0.00028610
         when "000101101010" => A <= "000000000001001000"; -- Line 2   Column 107   Coefficient 0.00027466
         when "000101101011" => A <= "000000000001000010"; -- Line 2   Column 108   Coefficient 0.00025177
         when "000101101100" => A <= "000000000001111110"; -- Line 2   Column 109   Coefficient 0.00048065
         when "000101101101" => A <= "000000000010010101"; -- Line 2   Column 110   Coefficient 0.00056839
         when "000101101110" => A <= "000000000001100101"; -- Line 2   Column 111   Coefficient 0.00038528
         when "000101101111" => A <= "000000000000110011"; -- Line 2   Column 112   Coefficient 0.00019455
         when "000101110000" => A <= "000000000000000111"; -- Line 2   Column 113   Coefficient 0.00002670
         when "000101110001" => A <= "111111111111100110"; -- Line 2   Column 114   Coefficient -0.00009918
         when "000101110010" => A <= "111111111111110100"; -- Line 2   Column 115   Coefficient -0.00004578
         when "000101110011" => A <= "000000000000000011"; -- Line 2   Column 116   Coefficient 0.00001144
         when "000101110100" => A <= "000000000000000100"; -- Line 2   Column 117   Coefficient 0.00001526
         when "000101110101" => A <= "000000000000000110"; -- Line 2   Column 118   Coefficient 0.00002289
         when "000101110110" => A <= "000000000000000011"; -- Line 2   Column 119   Coefficient 0.00001144
         when "000101110111" => A <= "111111111111111111"; -- Line 2   Column 120   Coefficient -0.00000381
         when "000101111000" => A <= "000000000000000000"; -- Line 2   Column 121   Coefficient 0.00000000
         when "000101111001" => A <= "000000000000000000"; -- Line 2   Column 122   Coefficient 0.00000000
         when "000101111010" => A <= "000000000000000000"; -- Line 2   Column 123   Coefficient 0.00000000
         when "000101111011" => A <= "000000000000000000"; -- Line 2   Column 124   Coefficient 0.00000000
         when "000101111100" => A <= "000000000000000000"; -- Line 2   Column 125   Coefficient 0.00000000
         when "000101111101" => A <= "000000000000000000"; -- Line 2   Column 126   Coefficient 0.00000000
         when "000101111110" => A <= "000000000000000000"; -- Line 2   Column 127   Coefficient 0.00000000
         when "000101111111" => A <= "000000000000000000"; -- Line 2   Column 128   Coefficient 0.00000000
         when "000110000000" => A <= "000000000000000000"; -- Line 2   Column 129   Coefficient 0.00000000
         when "000110000001" => A <= "000000000000000000"; -- Line 2   Column 130   Coefficient 0.00000000
         when "000110000010" => A <= "000000000000000000"; -- Line 2   Column 131   Coefficient 0.00000000
         when "000110000011" => A <= "000000000000000000"; -- Line 2   Column 132   Coefficient 0.00000000
         when "000110000100" => A <= "000000000000000000"; -- Line 2   Column 133   Coefficient 0.00000000
         when "000110000101" => A <= "000000000000000000"; -- Line 2   Column 134   Coefficient 0.00000000
         when "000110000110" => A <= "000000000000000000"; -- Line 2   Column 135   Coefficient 0.00000000
         when "000110000111" => A <= "000000000000000000"; -- Line 2   Column 136   Coefficient 0.00000000
         when "000110001000" => A <= "000000000000000000"; -- Line 2   Column 137   Coefficient 0.00000000
         when "000110001001" => A <= "000000000000000000"; -- Line 2   Column 138   Coefficient 0.00000000
         when "000110001010" => A <= "000000000000000000"; -- Line 2   Column 139   Coefficient 0.00000000
         when "000110001011" => A <= "000000000000000000"; -- Line 2   Column 140   Coefficient 0.00000000
         when "000110001100" => A <= "000000000000000000"; -- Line 2   Column 141   Coefficient 0.00000000
         when "000110001101" => A <= "000000000000000000"; -- Line 2   Column 142   Coefficient 0.00000000
         when "000110001110" => A <= "000000000000000000"; -- Line 2   Column 143   Coefficient 0.00000000
         when "000110001111" => A <= "000000000000000000"; -- Line 2   Column 144   Coefficient 0.00000000
         when "000110010000" => A <= "000000000000000000"; -- Line 2   Column 145   Coefficient 0.00000000
         when "000110010001" => A <= "000000000000000000"; -- Line 2   Column 146   Coefficient 0.00000000
         when "000110010010" => A <= "000000000000000000"; -- Line 2   Column 147   Coefficient 0.00000000
         when "000110010011" => A <= "000000000000000000"; -- Line 2   Column 148   Coefficient 0.00000000
         when "000110010100" => A <= "000000000000000000"; -- Line 2   Column 149   Coefficient 0.00000000
         when "000110010101" => A <= "000000000000000000"; -- Line 2   Column 150   Coefficient 0.00000000
         when "000110010110" => A <= "000000000000000000"; -- Line 2   Column 151   Coefficient 0.00000000
         when "000110010111" => A <= "000000000000000000"; -- Line 2   Column 152   Coefficient 0.00000000
         when "000110011000" => A <= "000000000000000000"; -- Line 2   Column 153   Coefficient 0.00000000
         when "000110011001" => A <= "000000000000000000"; -- Line 2   Column 154   Coefficient 0.00000000
         when "000110011010" => A <= "000000000000000000"; -- Line 2   Column 155   Coefficient 0.00000000
         when "000110011011" => A <= "000000000000000000"; -- Line 2   Column 156   Coefficient 0.00000000
         when "000110011100" => A <= "000000000000000000"; -- Line 2   Column 157   Coefficient 0.00000000
         when "000110011101" => A <= "000000000000000000"; -- Line 2   Column 158   Coefficient 0.00000000
         when "000110011110" => A <= "000000000000000000"; -- Line 2   Column 159   Coefficient 0.00000000
         when "000110011111" => A <= "000000000000000000"; -- Line 2   Column 160   Coefficient 0.00000000
         when "000110100000" => A <= "000000000000000000"; -- Line 2   Column 161   Coefficient 0.00000000
         when "000110100001" => A <= "000000000000000000"; -- Line 2   Column 162   Coefficient 0.00000000
         when "000110100010" => A <= "000000000000000000"; -- Line 2   Column 163   Coefficient 0.00000000
         when "000110100011" => A <= "000000000000000000"; -- Line 2   Column 164   Coefficient 0.00000000
         when "000110100100" => A <= "000000000000000000"; -- Line 2   Column 165   Coefficient 0.00000000
         when "000110100101" => A <= "000000000000000000"; -- Line 2   Column 166   Coefficient 0.00000000
         when "000110100110" => A <= "000000000000000000"; -- Line 2   Column 167   Coefficient 0.00000000
         when "000110100111" => A <= "000000000000000000"; -- Line 2   Column 168   Coefficient 0.00000000
         when "000110101000" => A <= "000000000000000000"; -- Line 2   Column 169   Coefficient 0.00000000
         when "000110101001" => A <= "000000000000000000"; -- Line 2   Column 170   Coefficient 0.00000000
         when "000110101010" => A <= "000000000000000000"; -- Line 2   Column 171   Coefficient 0.00000000
         when "000110101011" => A <= "000000000000000000"; -- Line 2   Column 172   Coefficient 0.00000000
         when "000110101100" => A <= "000000000000000000"; -- Line 2   Column 173   Coefficient 0.00000000
         when "000110101101" => A <= "000000000000000000"; -- Line 2   Column 174   Coefficient 0.00000000
         when "000110101110" => A <= "000000000000000000"; -- Line 2   Column 175   Coefficient 0.00000000
         when "000110101111" => A <= "000000000000000000"; -- Line 2   Column 176   Coefficient 0.00000000
         when "000110110000" => A <= "000000000000000000"; -- Line 2   Column 177   Coefficient 0.00000000
         when "000110110001" => A <= "000000000000000000"; -- Line 2   Column 178   Coefficient 0.00000000
         when "000110110010" => A <= "000000000000000000"; -- Line 2   Column 179   Coefficient 0.00000000
         when "000110110011" => A <= "000000000000000000"; -- Line 2   Column 180   Coefficient 0.00000000
         when "000110110100" => A <= "000000000000000000"; -- Line 2   Column 181   Coefficient 0.00000000
         when "000110110101" => A <= "000000000000000000"; -- Line 2   Column 182   Coefficient 0.00000000
         when "000110110110" => A <= "000000000000000000"; -- Line 2   Column 183   Coefficient 0.00000000
         when "000110110111" => A <= "000000000000000000"; -- Line 2   Column 184   Coefficient 0.00000000
         when "000110111000" => A <= "000000000000000000"; -- Line 2   Column 185   Coefficient 0.00000000
         when "000110111001" => A <= "000000000000000000"; -- Line 2   Column 186   Coefficient 0.00000000
         when "000110111010" => A <= "000000000000000000"; -- Line 2   Column 187   Coefficient 0.00000000
         when "000110111011" => A <= "000000000000000000"; -- Line 2   Column 188   Coefficient 0.00000000
         when "000110111100" => A <= "000000000000000000"; -- Line 2   Column 189   Coefficient 0.00000000
         when "000110111101" => A <= "000000000000000000"; -- Line 2   Column 190   Coefficient 0.00000000
         when "000110111110" => A <= "000000000000000000"; -- Line 2   Column 191   Coefficient 0.00000000
         when "000110111111" => A <= "000000000000000000"; -- Line 2   Column 192   Coefficient 0.00000000
         when "000111000000" => A <= "000000000000000000"; -- Line 2   Column 193   Coefficient 0.00000000
         when "000111000001" => A <= "000000000000000000"; -- Line 2   Column 194   Coefficient 0.00000000
         when "000111000010" => A <= "000000000000000000"; -- Line 2   Column 195   Coefficient 0.00000000
         when "000111000011" => A <= "000000000000000000"; -- Line 2   Column 196   Coefficient 0.00000000
         when "000111000100" => A <= "000000000000000000"; -- Line 2   Column 197   Coefficient 0.00000000
         when "000111000101" => A <= "000000000000000000"; -- Line 2   Column 198   Coefficient 0.00000000
         when "000111000110" => A <= "000000000000000000"; -- Line 2   Column 199   Coefficient 0.00000000
         when "000111000111" => A <= "000000000000000000"; -- Line 2   Column 200   Coefficient 0.00000000
         when "000111001000" => A <= "000000000000000000"; -- Line 2   Column 201   Coefficient 0.00000000
         when "000111001001" => A <= "000000000000000000"; -- Line 2   Column 202   Coefficient 0.00000000
         when "000111001010" => A <= "000000000000000000"; -- Line 2   Column 203   Coefficient 0.00000000
         when "000111001011" => A <= "000000000000000000"; -- Line 2   Column 204   Coefficient 0.00000000
         when "000111001100" => A <= "000000000000000000"; -- Line 2   Column 205   Coefficient 0.00000000
         when "000111001101" => A <= "000000000000000000"; -- Line 2   Column 206   Coefficient 0.00000000
         when "000111001110" => A <= "000000000000000000"; -- Line 2   Column 207   Coefficient 0.00000000
         when "000111001111" => A <= "000000000000000000"; -- Line 2   Column 208   Coefficient 0.00000000
         when "000111010000" => A <= "000000000000000000"; -- Line 2   Column 209   Coefficient 0.00000000
         when "000111010001" => A <= "000000000000000000"; -- Line 2   Column 210   Coefficient 0.00000000
         when "000111010010" => A <= "000000000000000000"; -- Line 2   Column 211   Coefficient 0.00000000
         when "000111010011" => A <= "000000000000000000"; -- Line 2   Column 212   Coefficient 0.00000000
         when "000111010100" => A <= "000000000000000000"; -- Line 2   Column 213   Coefficient 0.00000000
         when "000111010101" => A <= "000000000000000000"; -- Line 2   Column 214   Coefficient 0.00000000
         when "000111010110" => A <= "000000000000000000"; -- Line 2   Column 215   Coefficient 0.00000000
         when "000111010111" => A <= "000000000000000000"; -- Line 2   Column 216   Coefficient 0.00000000
         when "000111011000" => A <= "000000000000000000"; -- Line 2   Column 217   Coefficient 0.00000000
         when "000111011001" => A <= "000000000000000000"; -- Line 2   Column 218   Coefficient 0.00000000
         when "000111011010" => A <= "000000000000000000"; -- Line 2   Column 219   Coefficient 0.00000000
         when "000111011011" => A <= "000000000000000000"; -- Line 2   Column 220   Coefficient 0.00000000
         when "000111011100" => A <= "000000000000000000"; -- Line 2   Column 221   Coefficient 0.00000000
         when "000111011101" => A <= "000000000000000000"; -- Line 2   Column 222   Coefficient 0.00000000
         when "000111011110" => A <= "000000000000000000"; -- Line 2   Column 223   Coefficient 0.00000000
         when "000111011111" => A <= "000000000000000000"; -- Line 2   Column 224   Coefficient 0.00000000
         when "000111100000" => A <= "000000000000000000"; -- Line 2   Column 225   Coefficient 0.00000000
         when "000111100001" => A <= "000000000000000000"; -- Line 2   Column 226   Coefficient 0.00000000
         when "000111100010" => A <= "000000000000000000"; -- Line 2   Column 227   Coefficient 0.00000000
         when "000111100011" => A <= "000000000000000000"; -- Line 2   Column 228   Coefficient 0.00000000
         when "000111100100" => A <= "000000000000000000"; -- Line 2   Column 229   Coefficient 0.00000000
         when "000111100101" => A <= "000000000000000000"; -- Line 2   Column 230   Coefficient 0.00000000
         when "000111100110" => A <= "000000000000000000"; -- Line 2   Column 231   Coefficient 0.00000000
         when "000111100111" => A <= "000000000000000000"; -- Line 2   Column 232   Coefficient 0.00000000
         when "000111101000" => A <= "000000000000000000"; -- Line 2   Column 233   Coefficient 0.00000000
         when "000111101001" => A <= "000000000000000000"; -- Line 2   Column 234   Coefficient 0.00000000
         when "000111101010" => A <= "000000000000000000"; -- Line 2   Column 235   Coefficient 0.00000000
         when "000111101011" => A <= "000000000000000000"; -- Line 2   Column 236   Coefficient 0.00000000
         when "000111101100" => A <= "000000000000000000"; -- Line 2   Column 237   Coefficient 0.00000000
         when "000111101101" => A <= "000000000000000000"; -- Line 2   Column 238   Coefficient 0.00000000
         when "000111101110" => A <= "000000000000000000"; -- Line 2   Column 239   Coefficient 0.00000000
         when "000111101111" => A <= "000000000000000000"; -- Line 2   Column 240   Coefficient 0.00000000
         when "000111110000" => A <= "000000000000000000"; -- Line 2   Column 241   Coefficient 0.00000000
         when "000111110001" => A <= "000000000000000000"; -- Line 2   Column 242   Coefficient 0.00000000
         when "000111110010" => A <= "000000000000000000"; -- Line 2   Column 243   Coefficient 0.00000000
         when "000111110011" => A <= "000000000000000000"; -- Line 2   Column 244   Coefficient 0.00000000
         when "000111110100" => A <= "000000000000000000"; -- Line 2   Column 245   Coefficient 0.00000000
         when "000111110101" => A <= "000000000000000000"; -- Line 2   Column 246   Coefficient 0.00000000
         when "000111110110" => A <= "000000000000000000"; -- Line 2   Column 247   Coefficient 0.00000000
         when "000111110111" => A <= "000000000000000000"; -- Line 2   Column 248   Coefficient 0.00000000
         when "000111111000" => A <= "000000000000000000"; -- Line 2   Column 249   Coefficient 0.00000000
         when "000111111001" => A <= "000000000000000000"; -- Line 2   Column 250   Coefficient 0.00000000
         when "000111111010" => A <= "000000000000000000"; -- Line 2   Column 251   Coefficient 0.00000000
         when "000111111011" => A <= "000000000000000000"; -- Line 2   Column 252   Coefficient 0.00000000
         when "000111111100" => A <= "000000000000000000"; -- Line 2   Column 253   Coefficient 0.00000000
         when "000111111101" => A <= "000000000000000000"; -- Line 2   Column 254   Coefficient 0.00000000
         when "000111111110" => A <= "000000000000000000"; -- Line 2   Column 255   Coefficient 0.00000000
         when "000111111111" => A <= "000000000000000000"; -- Line 2   Column 256   Coefficient 0.00000000
         when "001000000000" => A <= "000000000000000000"; -- Line 3   Column 1   Coefficient 0.00000000
         when "001000000001" => A <= "000000000000000000"; -- Line 3   Column 2   Coefficient 0.00000000
         when "001000000010" => A <= "000000000000000000"; -- Line 3   Column 3   Coefficient 0.00000000
         when "001000000011" => A <= "000000000000000000"; -- Line 3   Column 4   Coefficient 0.00000000
         when "001000000100" => A <= "000000000000000000"; -- Line 3   Column 5   Coefficient 0.00000000
         when "001000000101" => A <= "000000000000000000"; -- Line 3   Column 6   Coefficient 0.00000000
         when "001000000110" => A <= "000000000000000000"; -- Line 3   Column 7   Coefficient 0.00000000
         when "001000000111" => A <= "000000000000000000"; -- Line 3   Column 8   Coefficient 0.00000000
         when "001000001000" => A <= "000000000000000000"; -- Line 3   Column 9   Coefficient 0.00000000
         when "001000001001" => A <= "000000000000000000"; -- Line 3   Column 10   Coefficient 0.00000000
         when "001000001010" => A <= "000000000000000000"; -- Line 3   Column 11   Coefficient 0.00000000
         when "001000001011" => A <= "000000000000000000"; -- Line 3   Column 12   Coefficient 0.00000000
         when "001000001100" => A <= "000000000000000000"; -- Line 3   Column 13   Coefficient 0.00000000
         when "001000001101" => A <= "000000000000000000"; -- Line 3   Column 14   Coefficient 0.00000000
         when "001000001110" => A <= "000000000000000000"; -- Line 3   Column 15   Coefficient 0.00000000
         when "001000001111" => A <= "000000000000000000"; -- Line 3   Column 16   Coefficient 0.00000000
         when "001000010000" => A <= "000000000000000000"; -- Line 3   Column 17   Coefficient 0.00000000
         when "001000010001" => A <= "000000000000000000"; -- Line 3   Column 18   Coefficient 0.00000000
         when "001000010010" => A <= "000000000000000000"; -- Line 3   Column 19   Coefficient 0.00000000
         when "001000010011" => A <= "000000000000000000"; -- Line 3   Column 20   Coefficient 0.00000000
         when "001000010100" => A <= "000000000000000000"; -- Line 3   Column 21   Coefficient 0.00000000
         when "001000010101" => A <= "000000000000000000"; -- Line 3   Column 22   Coefficient 0.00000000
         when "001000010110" => A <= "000000000000000000"; -- Line 3   Column 23   Coefficient 0.00000000
         when "001000010111" => A <= "000000000000000000"; -- Line 3   Column 24   Coefficient 0.00000000
         when "001000011000" => A <= "000000000000000000"; -- Line 3   Column 25   Coefficient 0.00000000
         when "001000011001" => A <= "000000000000000000"; -- Line 3   Column 26   Coefficient 0.00000000
         when "001000011010" => A <= "000000000000000000"; -- Line 3   Column 27   Coefficient 0.00000000
         when "001000011011" => A <= "000000000000000000"; -- Line 3   Column 28   Coefficient 0.00000000
         when "001000011100" => A <= "000000000000000000"; -- Line 3   Column 29   Coefficient 0.00000000
         when "001000011101" => A <= "000000000000000000"; -- Line 3   Column 30   Coefficient 0.00000000
         when "001000011110" => A <= "000000000000000000"; -- Line 3   Column 31   Coefficient 0.00000000
         when "001000011111" => A <= "000000000000000000"; -- Line 3   Column 32   Coefficient 0.00000000
         when "001000100000" => A <= "000000000000001001"; -- Line 3   Column 33   Coefficient 0.00003433
         when "001000100001" => A <= "000000000000000011"; -- Line 3   Column 34   Coefficient 0.00001144
         when "001000100010" => A <= "111111111111001011"; -- Line 3   Column 35   Coefficient -0.00020218
         when "001000100011" => A <= "111111111110100110"; -- Line 3   Column 36   Coefficient -0.00034332
         when "001000100100" => A <= "111111111110010010"; -- Line 3   Column 37   Coefficient -0.00041962
         when "001000100101" => A <= "111111111111010011"; -- Line 3   Column 38   Coefficient -0.00017166
         when "001000100110" => A <= "000000000011111000"; -- Line 3   Column 39   Coefficient 0.00094604
         when "001000100111" => A <= "000000001000010011"; -- Line 3   Column 40   Coefficient 0.00202560
         when "001000101000" => A <= "000000001010110110"; -- Line 3   Column 41   Coefficient 0.00264740
         when "001000101001" => A <= "000000001101001100"; -- Line 3   Column 42   Coefficient 0.00321960
         when "001000101010" => A <= "000000001111111100"; -- Line 3   Column 43   Coefficient 0.00389099
         when "001000101011" => A <= "000000010000011000"; -- Line 3   Column 44   Coefficient 0.00399780
         when "001000101100" => A <= "000000001111000010"; -- Line 3   Column 45   Coefficient 0.00366974
         when "001000101101" => A <= "000000000111011010"; -- Line 3   Column 46   Coefficient 0.00180817
         when "001000101110" => A <= "111111110001010101"; -- Line 3   Column 47   Coefficient -0.00358200
         when "001000101111" => A <= "111111011001111001"; -- Line 3   Column 48   Coefficient -0.00930405
         when "001000110000" => A <= "111111000100111001"; -- Line 3   Column 49   Coefficient -0.01443100
         when "001000110001" => A <= "111110110001100001"; -- Line 3   Column 50   Coefficient -0.01916122
         when "001000110010" => A <= "111110100110010011"; -- Line 3   Column 51   Coefficient -0.02190018
         when "001000110011" => A <= "111110011011111010"; -- Line 3   Column 52   Coefficient -0.02443695
         when "001000110100" => A <= "111110010000110000"; -- Line 3   Column 53   Coefficient -0.02716064
         when "001000110101" => A <= "111110000101010011"; -- Line 3   Column 54   Coefficient -0.02995682
         when "001000110110" => A <= "111101110100001010"; -- Line 3   Column 55   Coefficient -0.03414154
         when "001000110111" => A <= "111101100110110000"; -- Line 3   Column 56   Coefficient -0.03741455
         when "001000111000" => A <= "111101100010101111"; -- Line 3   Column 57   Coefficient -0.03839493
         when "001000111001" => A <= "111101100010001110"; -- Line 3   Column 58   Coefficient -0.03852081
         when "001000111010" => A <= "111101100000101101"; -- Line 3   Column 59   Coefficient -0.03889084
         when "001000111011" => A <= "111101101011101110"; -- Line 3   Column 60   Coefficient -0.03620148
         when "001000111100" => A <= "111110000010011110"; -- Line 3   Column 61   Coefficient -0.03064728
         when "001000111101" => A <= "111110110101100100"; -- Line 3   Column 62   Coefficient -0.01817322
         when "001000111110" => A <= "000000100101011001"; -- Line 3   Column 63   Coefficient 0.00912857
         when "001000111111" => A <= "000010011110111100"; -- Line 3   Column 64   Coefficient 0.03880310
         when "001001000000" => A <= "000100010010000101"; -- Line 3   Column 65   Coefficient 0.06691360
         when "001001000001" => A <= "000110000101110011"; -- Line 3   Column 66   Coefficient 0.09516525
         when "001001000010" => A <= "000111100110110001"; -- Line 3   Column 67   Coefficient 0.11883926
         when "001001000011" => A <= "001001000110101001"; -- Line 3   Column 68   Coefficient 0.14224625
         when "001001000100" => A <= "001010101100000111"; -- Line 3   Column 69   Coefficient 0.16701889
         when "001001000101" => A <= "001100001011101000"; -- Line 3   Column 70   Coefficient 0.19033813
         when "001001000110" => A <= "001101100011111111"; -- Line 3   Column 71   Coefficient 0.21191025
         when "001001000111" => A <= "001110110101010100"; -- Line 3   Column 72   Coefficient 0.23176575
         when "001001001000" => A <= "001111111010100001"; -- Line 3   Column 73   Coefficient 0.24866104
         when "001001001001" => A <= "010000111010100101"; -- Line 3   Column 74   Coefficient 0.26430130
         when "001001001010" => A <= "010010000001100011"; -- Line 3   Column 75   Coefficient 0.28162766
         when "001001001011" => A <= "010010110100110100"; -- Line 3   Column 76   Coefficient 0.29414368
         when "001001001100" => A <= "010011010010100110"; -- Line 3   Column 77   Coefficient 0.30141449
         when "001001001101" => A <= "010011000101100111"; -- Line 3   Column 78   Coefficient 0.29824448
         when "001001001110" => A <= "010001011110001011"; -- Line 3   Column 79   Coefficient 0.27299118
         when "001001001111" => A <= "001111100101110011"; -- Line 3   Column 80   Coefficient 0.24360275
         when "001001010000" => A <= "001101110100101001"; -- Line 3   Column 81   Coefficient 0.21597672
         when "001001010001" => A <= "001011111101111010"; -- Line 3   Column 82   Coefficient 0.18698883
         when "001001010010" => A <= "001010011001111000"; -- Line 3   Column 83   Coefficient 0.16256714
         when "001001010011" => A <= "001000110101000000"; -- Line 3   Column 84   Coefficient 0.13793945
         when "001001010100" => A <= "000111000101010101"; -- Line 3   Column 85   Coefficient 0.11067581
         when "001001010101" => A <= "000101100000010101"; -- Line 3   Column 86   Coefficient 0.08601761
         when "001001010110" => A <= "000100010011001101"; -- Line 3   Column 87   Coefficient 0.06718826
         when "001001010111" => A <= "000011001010010011"; -- Line 3   Column 88   Coefficient 0.04938889
         when "001001011000" => A <= "000010000100001011"; -- Line 3   Column 89   Coefficient 0.03226852
         when "001001011001" => A <= "000000111110100110"; -- Line 3   Column 90   Coefficient 0.01528168
         when "001001011010" => A <= "111111101010001000"; -- Line 3   Column 91   Coefficient -0.00534058
         when "001001011011" => A <= "111110100000101100"; -- Line 3   Column 92   Coefficient -0.02326965
         when "001001011100" => A <= "111101100111001110"; -- Line 3   Column 93   Coefficient -0.03730011
         when "001001011101" => A <= "111101000110110001"; -- Line 3   Column 94   Coefficient -0.04522324
         when "001001011110" => A <= "111101011101101101"; -- Line 3   Column 95   Coefficient -0.03962326
         when "001001011111" => A <= "111101111110110001"; -- Line 3   Column 96   Coefficient -0.03155136
         when "001001100000" => A <= "111110011010010101"; -- Line 3   Column 97   Coefficient -0.02482224
         when "001001100001" => A <= "111110111010000001"; -- Line 3   Column 98   Coefficient -0.01708603
         when "001001100010" => A <= "111111010000101110"; -- Line 3   Column 99   Coefficient -0.01154327
         when "001001100011" => A <= "111111100111100010"; -- Line 3   Column 100   Coefficient -0.00597382
         when "001001100100" => A <= "000000000100100100"; -- Line 3   Column 101   Coefficient 0.00111389
         when "001001100101" => A <= "000000011000110111"; -- Line 3   Column 102   Coefficient 0.00606918
         when "001001100110" => A <= "000000010111101010"; -- Line 3   Column 103   Coefficient 0.00577545
         when "001001100111" => A <= "000000010100111001"; -- Line 3   Column 104   Coefficient 0.00510025
         when "001001101000" => A <= "000000010100110111"; -- Line 3   Column 105   Coefficient 0.00509262
         when "001001101001" => A <= "000000010110010000"; -- Line 3   Column 106   Coefficient 0.00543213
         when "001001101010" => A <= "000000100010100100"; -- Line 3   Column 107   Coefficient 0.00843811
         when "001001101011" => A <= "000000101101010111"; -- Line 3   Column 108   Coefficient 0.01107407
         when "001001101100" => A <= "000000110010101110"; -- Line 3   Column 109   Coefficient 0.01238251
         when "001001101101" => A <= "000000110100010110"; -- Line 3   Column 110   Coefficient 0.01277924
         when "001001101110" => A <= "000000101011110101"; -- Line 3   Column 111   Coefficient 0.01070023
         when "001001101111" => A <= "000000100001110011"; -- Line 3   Column 112   Coefficient 0.00825119
         when "001001110000" => A <= "000000011001110100"; -- Line 3   Column 113   Coefficient 0.00630188
         when "001001110001" => A <= "000000010001001000"; -- Line 3   Column 114   Coefficient 0.00418091
         when "001001110010" => A <= "000000001001011000"; -- Line 3   Column 115   Coefficient 0.00228882
         when "001001110011" => A <= "000000000010010011"; -- Line 3   Column 116   Coefficient 0.00056076
         when "001001110100" => A <= "111111111010111001"; -- Line 3   Column 117   Coefficient -0.00124741
         when "001001110101" => A <= "111111110110011111"; -- Line 3   Column 118   Coefficient -0.00232315
         when "001001110110" => A <= "111111111001000110"; -- Line 3   Column 119   Coefficient -0.00168610
         when "001001110111" => A <= "111111111100011110"; -- Line 3   Column 120   Coefficient -0.00086212
         when "001001111000" => A <= "111111111110110111"; -- Line 3   Column 121   Coefficient -0.00027847
         when "001001111001" => A <= "000000000001001011"; -- Line 3   Column 122   Coefficient 0.00028610
         when "001001111010" => A <= "000000000001001000"; -- Line 3   Column 123   Coefficient 0.00027466
         when "001001111011" => A <= "000000000001000010"; -- Line 3   Column 124   Coefficient 0.00025177
         when "001001111100" => A <= "000000000001111110"; -- Line 3   Column 125   Coefficient 0.00048065
         when "001001111101" => A <= "000000000010010101"; -- Line 3   Column 126   Coefficient 0.00056839
         when "001001111110" => A <= "000000000001100101"; -- Line 3   Column 127   Coefficient 0.00038528
         when "001001111111" => A <= "000000000000110011"; -- Line 3   Column 128   Coefficient 0.00019455
         when "001010000000" => A <= "000000000000000111"; -- Line 3   Column 129   Coefficient 0.00002670
         when "001010000001" => A <= "111111111111100110"; -- Line 3   Column 130   Coefficient -0.00009918
         when "001010000010" => A <= "111111111111110100"; -- Line 3   Column 131   Coefficient -0.00004578
         when "001010000011" => A <= "000000000000000011"; -- Line 3   Column 132   Coefficient 0.00001144
         when "001010000100" => A <= "000000000000000100"; -- Line 3   Column 133   Coefficient 0.00001526
         when "001010000101" => A <= "000000000000000110"; -- Line 3   Column 134   Coefficient 0.00002289
         when "001010000110" => A <= "000000000000000011"; -- Line 3   Column 135   Coefficient 0.00001144
         when "001010000111" => A <= "111111111111111111"; -- Line 3   Column 136   Coefficient -0.00000381
         when "001010001000" => A <= "000000000000000000"; -- Line 3   Column 137   Coefficient 0.00000000
         when "001010001001" => A <= "000000000000000000"; -- Line 3   Column 138   Coefficient 0.00000000
         when "001010001010" => A <= "000000000000000000"; -- Line 3   Column 139   Coefficient 0.00000000
         when "001010001011" => A <= "000000000000000000"; -- Line 3   Column 140   Coefficient 0.00000000
         when "001010001100" => A <= "000000000000000000"; -- Line 3   Column 141   Coefficient 0.00000000
         when "001010001101" => A <= "000000000000000000"; -- Line 3   Column 142   Coefficient 0.00000000
         when "001010001110" => A <= "000000000000000000"; -- Line 3   Column 143   Coefficient 0.00000000
         when "001010001111" => A <= "000000000000000000"; -- Line 3   Column 144   Coefficient 0.00000000
         when "001010010000" => A <= "000000000000000000"; -- Line 3   Column 145   Coefficient 0.00000000
         when "001010010001" => A <= "000000000000000000"; -- Line 3   Column 146   Coefficient 0.00000000
         when "001010010010" => A <= "000000000000000000"; -- Line 3   Column 147   Coefficient 0.00000000
         when "001010010011" => A <= "000000000000000000"; -- Line 3   Column 148   Coefficient 0.00000000
         when "001010010100" => A <= "000000000000000000"; -- Line 3   Column 149   Coefficient 0.00000000
         when "001010010101" => A <= "000000000000000000"; -- Line 3   Column 150   Coefficient 0.00000000
         when "001010010110" => A <= "000000000000000000"; -- Line 3   Column 151   Coefficient 0.00000000
         when "001010010111" => A <= "000000000000000000"; -- Line 3   Column 152   Coefficient 0.00000000
         when "001010011000" => A <= "000000000000000000"; -- Line 3   Column 153   Coefficient 0.00000000
         when "001010011001" => A <= "000000000000000000"; -- Line 3   Column 154   Coefficient 0.00000000
         when "001010011010" => A <= "000000000000000000"; -- Line 3   Column 155   Coefficient 0.00000000
         when "001010011011" => A <= "000000000000000000"; -- Line 3   Column 156   Coefficient 0.00000000
         when "001010011100" => A <= "000000000000000000"; -- Line 3   Column 157   Coefficient 0.00000000
         when "001010011101" => A <= "000000000000000000"; -- Line 3   Column 158   Coefficient 0.00000000
         when "001010011110" => A <= "000000000000000000"; -- Line 3   Column 159   Coefficient 0.00000000
         when "001010011111" => A <= "000000000000000000"; -- Line 3   Column 160   Coefficient 0.00000000
         when "001010100000" => A <= "000000000000000000"; -- Line 3   Column 161   Coefficient 0.00000000
         when "001010100001" => A <= "000000000000000000"; -- Line 3   Column 162   Coefficient 0.00000000
         when "001010100010" => A <= "000000000000000000"; -- Line 3   Column 163   Coefficient 0.00000000
         when "001010100011" => A <= "000000000000000000"; -- Line 3   Column 164   Coefficient 0.00000000
         when "001010100100" => A <= "000000000000000000"; -- Line 3   Column 165   Coefficient 0.00000000
         when "001010100101" => A <= "000000000000000000"; -- Line 3   Column 166   Coefficient 0.00000000
         when "001010100110" => A <= "000000000000000000"; -- Line 3   Column 167   Coefficient 0.00000000
         when "001010100111" => A <= "000000000000000000"; -- Line 3   Column 168   Coefficient 0.00000000
         when "001010101000" => A <= "000000000000000000"; -- Line 3   Column 169   Coefficient 0.00000000
         when "001010101001" => A <= "000000000000000000"; -- Line 3   Column 170   Coefficient 0.00000000
         when "001010101010" => A <= "000000000000000000"; -- Line 3   Column 171   Coefficient 0.00000000
         when "001010101011" => A <= "000000000000000000"; -- Line 3   Column 172   Coefficient 0.00000000
         when "001010101100" => A <= "000000000000000000"; -- Line 3   Column 173   Coefficient 0.00000000
         when "001010101101" => A <= "000000000000000000"; -- Line 3   Column 174   Coefficient 0.00000000
         when "001010101110" => A <= "000000000000000000"; -- Line 3   Column 175   Coefficient 0.00000000
         when "001010101111" => A <= "000000000000000000"; -- Line 3   Column 176   Coefficient 0.00000000
         when "001010110000" => A <= "000000000000000000"; -- Line 3   Column 177   Coefficient 0.00000000
         when "001010110001" => A <= "000000000000000000"; -- Line 3   Column 178   Coefficient 0.00000000
         when "001010110010" => A <= "000000000000000000"; -- Line 3   Column 179   Coefficient 0.00000000
         when "001010110011" => A <= "000000000000000000"; -- Line 3   Column 180   Coefficient 0.00000000
         when "001010110100" => A <= "000000000000000000"; -- Line 3   Column 181   Coefficient 0.00000000
         when "001010110101" => A <= "000000000000000000"; -- Line 3   Column 182   Coefficient 0.00000000
         when "001010110110" => A <= "000000000000000000"; -- Line 3   Column 183   Coefficient 0.00000000
         when "001010110111" => A <= "000000000000000000"; -- Line 3   Column 184   Coefficient 0.00000000
         when "001010111000" => A <= "000000000000000000"; -- Line 3   Column 185   Coefficient 0.00000000
         when "001010111001" => A <= "000000000000000000"; -- Line 3   Column 186   Coefficient 0.00000000
         when "001010111010" => A <= "000000000000000000"; -- Line 3   Column 187   Coefficient 0.00000000
         when "001010111011" => A <= "000000000000000000"; -- Line 3   Column 188   Coefficient 0.00000000
         when "001010111100" => A <= "000000000000000000"; -- Line 3   Column 189   Coefficient 0.00000000
         when "001010111101" => A <= "000000000000000000"; -- Line 3   Column 190   Coefficient 0.00000000
         when "001010111110" => A <= "000000000000000000"; -- Line 3   Column 191   Coefficient 0.00000000
         when "001010111111" => A <= "000000000000000000"; -- Line 3   Column 192   Coefficient 0.00000000
         when "001011000000" => A <= "000000000000000000"; -- Line 3   Column 193   Coefficient 0.00000000
         when "001011000001" => A <= "000000000000000000"; -- Line 3   Column 194   Coefficient 0.00000000
         when "001011000010" => A <= "000000000000000000"; -- Line 3   Column 195   Coefficient 0.00000000
         when "001011000011" => A <= "000000000000000000"; -- Line 3   Column 196   Coefficient 0.00000000
         when "001011000100" => A <= "000000000000000000"; -- Line 3   Column 197   Coefficient 0.00000000
         when "001011000101" => A <= "000000000000000000"; -- Line 3   Column 198   Coefficient 0.00000000
         when "001011000110" => A <= "000000000000000000"; -- Line 3   Column 199   Coefficient 0.00000000
         when "001011000111" => A <= "000000000000000000"; -- Line 3   Column 200   Coefficient 0.00000000
         when "001011001000" => A <= "000000000000000000"; -- Line 3   Column 201   Coefficient 0.00000000
         when "001011001001" => A <= "000000000000000000"; -- Line 3   Column 202   Coefficient 0.00000000
         when "001011001010" => A <= "000000000000000000"; -- Line 3   Column 203   Coefficient 0.00000000
         when "001011001011" => A <= "000000000000000000"; -- Line 3   Column 204   Coefficient 0.00000000
         when "001011001100" => A <= "000000000000000000"; -- Line 3   Column 205   Coefficient 0.00000000
         when "001011001101" => A <= "000000000000000000"; -- Line 3   Column 206   Coefficient 0.00000000
         when "001011001110" => A <= "000000000000000000"; -- Line 3   Column 207   Coefficient 0.00000000
         when "001011001111" => A <= "000000000000000000"; -- Line 3   Column 208   Coefficient 0.00000000
         when "001011010000" => A <= "000000000000000000"; -- Line 3   Column 209   Coefficient 0.00000000
         when "001011010001" => A <= "000000000000000000"; -- Line 3   Column 210   Coefficient 0.00000000
         when "001011010010" => A <= "000000000000000000"; -- Line 3   Column 211   Coefficient 0.00000000
         when "001011010011" => A <= "000000000000000000"; -- Line 3   Column 212   Coefficient 0.00000000
         when "001011010100" => A <= "000000000000000000"; -- Line 3   Column 213   Coefficient 0.00000000
         when "001011010101" => A <= "000000000000000000"; -- Line 3   Column 214   Coefficient 0.00000000
         when "001011010110" => A <= "000000000000000000"; -- Line 3   Column 215   Coefficient 0.00000000
         when "001011010111" => A <= "000000000000000000"; -- Line 3   Column 216   Coefficient 0.00000000
         when "001011011000" => A <= "000000000000000000"; -- Line 3   Column 217   Coefficient 0.00000000
         when "001011011001" => A <= "000000000000000000"; -- Line 3   Column 218   Coefficient 0.00000000
         when "001011011010" => A <= "000000000000000000"; -- Line 3   Column 219   Coefficient 0.00000000
         when "001011011011" => A <= "000000000000000000"; -- Line 3   Column 220   Coefficient 0.00000000
         when "001011011100" => A <= "000000000000000000"; -- Line 3   Column 221   Coefficient 0.00000000
         when "001011011101" => A <= "000000000000000000"; -- Line 3   Column 222   Coefficient 0.00000000
         when "001011011110" => A <= "000000000000000000"; -- Line 3   Column 223   Coefficient 0.00000000
         when "001011011111" => A <= "000000000000000000"; -- Line 3   Column 224   Coefficient 0.00000000
         when "001011100000" => A <= "000000000000000000"; -- Line 3   Column 225   Coefficient 0.00000000
         when "001011100001" => A <= "000000000000000000"; -- Line 3   Column 226   Coefficient 0.00000000
         when "001011100010" => A <= "000000000000000000"; -- Line 3   Column 227   Coefficient 0.00000000
         when "001011100011" => A <= "000000000000000000"; -- Line 3   Column 228   Coefficient 0.00000000
         when "001011100100" => A <= "000000000000000000"; -- Line 3   Column 229   Coefficient 0.00000000
         when "001011100101" => A <= "000000000000000000"; -- Line 3   Column 230   Coefficient 0.00000000
         when "001011100110" => A <= "000000000000000000"; -- Line 3   Column 231   Coefficient 0.00000000
         when "001011100111" => A <= "000000000000000000"; -- Line 3   Column 232   Coefficient 0.00000000
         when "001011101000" => A <= "000000000000000000"; -- Line 3   Column 233   Coefficient 0.00000000
         when "001011101001" => A <= "000000000000000000"; -- Line 3   Column 234   Coefficient 0.00000000
         when "001011101010" => A <= "000000000000000000"; -- Line 3   Column 235   Coefficient 0.00000000
         when "001011101011" => A <= "000000000000000000"; -- Line 3   Column 236   Coefficient 0.00000000
         when "001011101100" => A <= "000000000000000000"; -- Line 3   Column 237   Coefficient 0.00000000
         when "001011101101" => A <= "000000000000000000"; -- Line 3   Column 238   Coefficient 0.00000000
         when "001011101110" => A <= "000000000000000000"; -- Line 3   Column 239   Coefficient 0.00000000
         when "001011101111" => A <= "000000000000000000"; -- Line 3   Column 240   Coefficient 0.00000000
         when "001011110000" => A <= "000000000000000000"; -- Line 3   Column 241   Coefficient 0.00000000
         when "001011110001" => A <= "000000000000000000"; -- Line 3   Column 242   Coefficient 0.00000000
         when "001011110010" => A <= "000000000000000000"; -- Line 3   Column 243   Coefficient 0.00000000
         when "001011110011" => A <= "000000000000000000"; -- Line 3   Column 244   Coefficient 0.00000000
         when "001011110100" => A <= "000000000000000000"; -- Line 3   Column 245   Coefficient 0.00000000
         when "001011110101" => A <= "000000000000000000"; -- Line 3   Column 246   Coefficient 0.00000000
         when "001011110110" => A <= "000000000000000000"; -- Line 3   Column 247   Coefficient 0.00000000
         when "001011110111" => A <= "000000000000000000"; -- Line 3   Column 248   Coefficient 0.00000000
         when "001011111000" => A <= "000000000000000000"; -- Line 3   Column 249   Coefficient 0.00000000
         when "001011111001" => A <= "000000000000000000"; -- Line 3   Column 250   Coefficient 0.00000000
         when "001011111010" => A <= "000000000000000000"; -- Line 3   Column 251   Coefficient 0.00000000
         when "001011111011" => A <= "000000000000000000"; -- Line 3   Column 252   Coefficient 0.00000000
         when "001011111100" => A <= "000000000000000000"; -- Line 3   Column 253   Coefficient 0.00000000
         when "001011111101" => A <= "000000000000000000"; -- Line 3   Column 254   Coefficient 0.00000000
         when "001011111110" => A <= "000000000000000000"; -- Line 3   Column 255   Coefficient 0.00000000
         when "001011111111" => A <= "000000000000000000"; -- Line 3   Column 256   Coefficient 0.00000000
         when "001100000000" => A <= "000000000000000000"; -- Line 4   Column 1   Coefficient 0.00000000
         when "001100000001" => A <= "000000000000000000"; -- Line 4   Column 2   Coefficient 0.00000000
         when "001100000010" => A <= "000000000000000000"; -- Line 4   Column 3   Coefficient 0.00000000
         when "001100000011" => A <= "000000000000000000"; -- Line 4   Column 4   Coefficient 0.00000000
         when "001100000100" => A <= "000000000000000000"; -- Line 4   Column 5   Coefficient 0.00000000
         when "001100000101" => A <= "000000000000000000"; -- Line 4   Column 6   Coefficient 0.00000000
         when "001100000110" => A <= "000000000000000000"; -- Line 4   Column 7   Coefficient 0.00000000
         when "001100000111" => A <= "000000000000000000"; -- Line 4   Column 8   Coefficient 0.00000000
         when "001100001000" => A <= "000000000000000000"; -- Line 4   Column 9   Coefficient 0.00000000
         when "001100001001" => A <= "000000000000000000"; -- Line 4   Column 10   Coefficient 0.00000000
         when "001100001010" => A <= "000000000000000000"; -- Line 4   Column 11   Coefficient 0.00000000
         when "001100001011" => A <= "000000000000000000"; -- Line 4   Column 12   Coefficient 0.00000000
         when "001100001100" => A <= "000000000000000000"; -- Line 4   Column 13   Coefficient 0.00000000
         when "001100001101" => A <= "000000000000000000"; -- Line 4   Column 14   Coefficient 0.00000000
         when "001100001110" => A <= "000000000000000000"; -- Line 4   Column 15   Coefficient 0.00000000
         when "001100001111" => A <= "000000000000000000"; -- Line 4   Column 16   Coefficient 0.00000000
         when "001100010000" => A <= "000000000000000000"; -- Line 4   Column 17   Coefficient 0.00000000
         when "001100010001" => A <= "000000000000000000"; -- Line 4   Column 18   Coefficient 0.00000000
         when "001100010010" => A <= "000000000000000000"; -- Line 4   Column 19   Coefficient 0.00000000
         when "001100010011" => A <= "000000000000000000"; -- Line 4   Column 20   Coefficient 0.00000000
         when "001100010100" => A <= "000000000000000000"; -- Line 4   Column 21   Coefficient 0.00000000
         when "001100010101" => A <= "000000000000000000"; -- Line 4   Column 22   Coefficient 0.00000000
         when "001100010110" => A <= "000000000000000000"; -- Line 4   Column 23   Coefficient 0.00000000
         when "001100010111" => A <= "000000000000000000"; -- Line 4   Column 24   Coefficient 0.00000000
         when "001100011000" => A <= "000000000000000000"; -- Line 4   Column 25   Coefficient 0.00000000
         when "001100011001" => A <= "000000000000000000"; -- Line 4   Column 26   Coefficient 0.00000000
         when "001100011010" => A <= "000000000000000000"; -- Line 4   Column 27   Coefficient 0.00000000
         when "001100011011" => A <= "000000000000000000"; -- Line 4   Column 28   Coefficient 0.00000000
         when "001100011100" => A <= "000000000000000000"; -- Line 4   Column 29   Coefficient 0.00000000
         when "001100011101" => A <= "000000000000000000"; -- Line 4   Column 30   Coefficient 0.00000000
         when "001100011110" => A <= "000000000000000000"; -- Line 4   Column 31   Coefficient 0.00000000
         when "001100011111" => A <= "000000000000000000"; -- Line 4   Column 32   Coefficient 0.00000000
         when "001100100000" => A <= "000000000000000000"; -- Line 4   Column 33   Coefficient 0.00000000
         when "001100100001" => A <= "000000000000000000"; -- Line 4   Column 34   Coefficient 0.00000000
         when "001100100010" => A <= "000000000000000000"; -- Line 4   Column 35   Coefficient 0.00000000
         when "001100100011" => A <= "000000000000000000"; -- Line 4   Column 36   Coefficient 0.00000000
         when "001100100100" => A <= "000000000000000000"; -- Line 4   Column 37   Coefficient 0.00000000
         when "001100100101" => A <= "000000000000000000"; -- Line 4   Column 38   Coefficient 0.00000000
         when "001100100110" => A <= "000000000000000000"; -- Line 4   Column 39   Coefficient 0.00000000
         when "001100100111" => A <= "000000000000000000"; -- Line 4   Column 40   Coefficient 0.00000000
         when "001100101000" => A <= "000000000000000000"; -- Line 4   Column 41   Coefficient 0.00000000
         when "001100101001" => A <= "000000000000000000"; -- Line 4   Column 42   Coefficient 0.00000000
         when "001100101010" => A <= "000000000000000000"; -- Line 4   Column 43   Coefficient 0.00000000
         when "001100101011" => A <= "000000000000000000"; -- Line 4   Column 44   Coefficient 0.00000000
         when "001100101100" => A <= "000000000000000000"; -- Line 4   Column 45   Coefficient 0.00000000
         when "001100101101" => A <= "000000000000000000"; -- Line 4   Column 46   Coefficient 0.00000000
         when "001100101110" => A <= "000000000000000000"; -- Line 4   Column 47   Coefficient 0.00000000
         when "001100101111" => A <= "000000000000000000"; -- Line 4   Column 48   Coefficient 0.00000000
         when "001100110000" => A <= "000000000000001001"; -- Line 4   Column 49   Coefficient 0.00003433
         when "001100110001" => A <= "000000000000000011"; -- Line 4   Column 50   Coefficient 0.00001144
         when "001100110010" => A <= "111111111111001011"; -- Line 4   Column 51   Coefficient -0.00020218
         when "001100110011" => A <= "111111111110100110"; -- Line 4   Column 52   Coefficient -0.00034332
         when "001100110100" => A <= "111111111110010010"; -- Line 4   Column 53   Coefficient -0.00041962
         when "001100110101" => A <= "111111111111010011"; -- Line 4   Column 54   Coefficient -0.00017166
         when "001100110110" => A <= "000000000011111000"; -- Line 4   Column 55   Coefficient 0.00094604
         when "001100110111" => A <= "000000001000010011"; -- Line 4   Column 56   Coefficient 0.00202560
         when "001100111000" => A <= "000000001010110110"; -- Line 4   Column 57   Coefficient 0.00264740
         when "001100111001" => A <= "000000001101001100"; -- Line 4   Column 58   Coefficient 0.00321960
         when "001100111010" => A <= "000000001111111100"; -- Line 4   Column 59   Coefficient 0.00389099
         when "001100111011" => A <= "000000010000011000"; -- Line 4   Column 60   Coefficient 0.00399780
         when "001100111100" => A <= "000000001111000010"; -- Line 4   Column 61   Coefficient 0.00366974
         when "001100111101" => A <= "000000000111011010"; -- Line 4   Column 62   Coefficient 0.00180817
         when "001100111110" => A <= "111111110001010101"; -- Line 4   Column 63   Coefficient -0.00358200
         when "001100111111" => A <= "111111011001111001"; -- Line 4   Column 64   Coefficient -0.00930405
         when "001101000000" => A <= "111111000100111001"; -- Line 4   Column 65   Coefficient -0.01443100
         when "001101000001" => A <= "111110110001100001"; -- Line 4   Column 66   Coefficient -0.01916122
         when "001101000010" => A <= "111110100110010011"; -- Line 4   Column 67   Coefficient -0.02190018
         when "001101000011" => A <= "111110011011111010"; -- Line 4   Column 68   Coefficient -0.02443695
         when "001101000100" => A <= "111110010000110000"; -- Line 4   Column 69   Coefficient -0.02716064
         when "001101000101" => A <= "111110000101010011"; -- Line 4   Column 70   Coefficient -0.02995682
         when "001101000110" => A <= "111101110100001010"; -- Line 4   Column 71   Coefficient -0.03414154
         when "001101000111" => A <= "111101100110110000"; -- Line 4   Column 72   Coefficient -0.03741455
         when "001101001000" => A <= "111101100010101111"; -- Line 4   Column 73   Coefficient -0.03839493
         when "001101001001" => A <= "111101100010001110"; -- Line 4   Column 74   Coefficient -0.03852081
         when "001101001010" => A <= "111101100000101101"; -- Line 4   Column 75   Coefficient -0.03889084
         when "001101001011" => A <= "111101101011101110"; -- Line 4   Column 76   Coefficient -0.03620148
         when "001101001100" => A <= "111110000010011110"; -- Line 4   Column 77   Coefficient -0.03064728
         when "001101001101" => A <= "111110110101100100"; -- Line 4   Column 78   Coefficient -0.01817322
         when "001101001110" => A <= "000000100101011001"; -- Line 4   Column 79   Coefficient 0.00912857
         when "001101001111" => A <= "000010011110111100"; -- Line 4   Column 80   Coefficient 0.03880310
         when "001101010000" => A <= "000100010010000101"; -- Line 4   Column 81   Coefficient 0.06691360
         when "001101010001" => A <= "000110000101110011"; -- Line 4   Column 82   Coefficient 0.09516525
         when "001101010010" => A <= "000111100110110001"; -- Line 4   Column 83   Coefficient 0.11883926
         when "001101010011" => A <= "001001000110101001"; -- Line 4   Column 84   Coefficient 0.14224625
         when "001101010100" => A <= "001010101100000111"; -- Line 4   Column 85   Coefficient 0.16701889
         when "001101010101" => A <= "001100001011101000"; -- Line 4   Column 86   Coefficient 0.19033813
         when "001101010110" => A <= "001101100011111111"; -- Line 4   Column 87   Coefficient 0.21191025
         when "001101010111" => A <= "001110110101010100"; -- Line 4   Column 88   Coefficient 0.23176575
         when "001101011000" => A <= "001111111010100001"; -- Line 4   Column 89   Coefficient 0.24866104
         when "001101011001" => A <= "010000111010100101"; -- Line 4   Column 90   Coefficient 0.26430130
         when "001101011010" => A <= "010010000001100011"; -- Line 4   Column 91   Coefficient 0.28162766
         when "001101011011" => A <= "010010110100110100"; -- Line 4   Column 92   Coefficient 0.29414368
         when "001101011100" => A <= "010011010010100110"; -- Line 4   Column 93   Coefficient 0.30141449
         when "001101011101" => A <= "010011000101100111"; -- Line 4   Column 94   Coefficient 0.29824448
         when "001101011110" => A <= "010001011110001011"; -- Line 4   Column 95   Coefficient 0.27299118
         when "001101011111" => A <= "001111100101110011"; -- Line 4   Column 96   Coefficient 0.24360275
         when "001101100000" => A <= "001101110100101001"; -- Line 4   Column 97   Coefficient 0.21597672
         when "001101100001" => A <= "001011111101111010"; -- Line 4   Column 98   Coefficient 0.18698883
         when "001101100010" => A <= "001010011001111000"; -- Line 4   Column 99   Coefficient 0.16256714
         when "001101100011" => A <= "001000110101000000"; -- Line 4   Column 100   Coefficient 0.13793945
         when "001101100100" => A <= "000111000101010101"; -- Line 4   Column 101   Coefficient 0.11067581
         when "001101100101" => A <= "000101100000010101"; -- Line 4   Column 102   Coefficient 0.08601761
         when "001101100110" => A <= "000100010011001101"; -- Line 4   Column 103   Coefficient 0.06718826
         when "001101100111" => A <= "000011001010010011"; -- Line 4   Column 104   Coefficient 0.04938889
         when "001101101000" => A <= "000010000100001011"; -- Line 4   Column 105   Coefficient 0.03226852
         when "001101101001" => A <= "000000111110100110"; -- Line 4   Column 106   Coefficient 0.01528168
         when "001101101010" => A <= "111111101010001000"; -- Line 4   Column 107   Coefficient -0.00534058
         when "001101101011" => A <= "111110100000101100"; -- Line 4   Column 108   Coefficient -0.02326965
         when "001101101100" => A <= "111101100111001110"; -- Line 4   Column 109   Coefficient -0.03730011
         when "001101101101" => A <= "111101000110110001"; -- Line 4   Column 110   Coefficient -0.04522324
         when "001101101110" => A <= "111101011101101101"; -- Line 4   Column 111   Coefficient -0.03962326
         when "001101101111" => A <= "111101111110110001"; -- Line 4   Column 112   Coefficient -0.03155136
         when "001101110000" => A <= "111110011010010101"; -- Line 4   Column 113   Coefficient -0.02482224
         when "001101110001" => A <= "111110111010000001"; -- Line 4   Column 114   Coefficient -0.01708603
         when "001101110010" => A <= "111111010000101110"; -- Line 4   Column 115   Coefficient -0.01154327
         when "001101110011" => A <= "111111100111100010"; -- Line 4   Column 116   Coefficient -0.00597382
         when "001101110100" => A <= "000000000100100100"; -- Line 4   Column 117   Coefficient 0.00111389
         when "001101110101" => A <= "000000011000110111"; -- Line 4   Column 118   Coefficient 0.00606918
         when "001101110110" => A <= "000000010111101010"; -- Line 4   Column 119   Coefficient 0.00577545
         when "001101110111" => A <= "000000010100111001"; -- Line 4   Column 120   Coefficient 0.00510025
         when "001101111000" => A <= "000000010100110111"; -- Line 4   Column 121   Coefficient 0.00509262
         when "001101111001" => A <= "000000010110010000"; -- Line 4   Column 122   Coefficient 0.00543213
         when "001101111010" => A <= "000000100010100100"; -- Line 4   Column 123   Coefficient 0.00843811
         when "001101111011" => A <= "000000101101010111"; -- Line 4   Column 124   Coefficient 0.01107407
         when "001101111100" => A <= "000000110010101110"; -- Line 4   Column 125   Coefficient 0.01238251
         when "001101111101" => A <= "000000110100010110"; -- Line 4   Column 126   Coefficient 0.01277924
         when "001101111110" => A <= "000000101011110101"; -- Line 4   Column 127   Coefficient 0.01070023
         when "001101111111" => A <= "000000100001110011"; -- Line 4   Column 128   Coefficient 0.00825119
         when "001110000000" => A <= "000000011001110100"; -- Line 4   Column 129   Coefficient 0.00630188
         when "001110000001" => A <= "000000010001001000"; -- Line 4   Column 130   Coefficient 0.00418091
         when "001110000010" => A <= "000000001001011000"; -- Line 4   Column 131   Coefficient 0.00228882
         when "001110000011" => A <= "000000000010010011"; -- Line 4   Column 132   Coefficient 0.00056076
         when "001110000100" => A <= "111111111010111001"; -- Line 4   Column 133   Coefficient -0.00124741
         when "001110000101" => A <= "111111110110011111"; -- Line 4   Column 134   Coefficient -0.00232315
         when "001110000110" => A <= "111111111001000110"; -- Line 4   Column 135   Coefficient -0.00168610
         when "001110000111" => A <= "111111111100011110"; -- Line 4   Column 136   Coefficient -0.00086212
         when "001110001000" => A <= "111111111110110111"; -- Line 4   Column 137   Coefficient -0.00027847
         when "001110001001" => A <= "000000000001001011"; -- Line 4   Column 138   Coefficient 0.00028610
         when "001110001010" => A <= "000000000001001000"; -- Line 4   Column 139   Coefficient 0.00027466
         when "001110001011" => A <= "000000000001000010"; -- Line 4   Column 140   Coefficient 0.00025177
         when "001110001100" => A <= "000000000001111110"; -- Line 4   Column 141   Coefficient 0.00048065
         when "001110001101" => A <= "000000000010010101"; -- Line 4   Column 142   Coefficient 0.00056839
         when "001110001110" => A <= "000000000001100101"; -- Line 4   Column 143   Coefficient 0.00038528
         when "001110001111" => A <= "000000000000110011"; -- Line 4   Column 144   Coefficient 0.00019455
         when "001110010000" => A <= "000000000000000111"; -- Line 4   Column 145   Coefficient 0.00002670
         when "001110010001" => A <= "111111111111100110"; -- Line 4   Column 146   Coefficient -0.00009918
         when "001110010010" => A <= "111111111111110100"; -- Line 4   Column 147   Coefficient -0.00004578
         when "001110010011" => A <= "000000000000000011"; -- Line 4   Column 148   Coefficient 0.00001144
         when "001110010100" => A <= "000000000000000100"; -- Line 4   Column 149   Coefficient 0.00001526
         when "001110010101" => A <= "000000000000000110"; -- Line 4   Column 150   Coefficient 0.00002289
         when "001110010110" => A <= "000000000000000011"; -- Line 4   Column 151   Coefficient 0.00001144
         when "001110010111" => A <= "111111111111111111"; -- Line 4   Column 152   Coefficient -0.00000381
         when "001110011000" => A <= "000000000000000000"; -- Line 4   Column 153   Coefficient 0.00000000
         when "001110011001" => A <= "000000000000000000"; -- Line 4   Column 154   Coefficient 0.00000000
         when "001110011010" => A <= "000000000000000000"; -- Line 4   Column 155   Coefficient 0.00000000
         when "001110011011" => A <= "000000000000000000"; -- Line 4   Column 156   Coefficient 0.00000000
         when "001110011100" => A <= "000000000000000000"; -- Line 4   Column 157   Coefficient 0.00000000
         when "001110011101" => A <= "000000000000000000"; -- Line 4   Column 158   Coefficient 0.00000000
         when "001110011110" => A <= "000000000000000000"; -- Line 4   Column 159   Coefficient 0.00000000
         when "001110011111" => A <= "000000000000000000"; -- Line 4   Column 160   Coefficient 0.00000000
         when "001110100000" => A <= "000000000000000000"; -- Line 4   Column 161   Coefficient 0.00000000
         when "001110100001" => A <= "000000000000000000"; -- Line 4   Column 162   Coefficient 0.00000000
         when "001110100010" => A <= "000000000000000000"; -- Line 4   Column 163   Coefficient 0.00000000
         when "001110100011" => A <= "000000000000000000"; -- Line 4   Column 164   Coefficient 0.00000000
         when "001110100100" => A <= "000000000000000000"; -- Line 4   Column 165   Coefficient 0.00000000
         when "001110100101" => A <= "000000000000000000"; -- Line 4   Column 166   Coefficient 0.00000000
         when "001110100110" => A <= "000000000000000000"; -- Line 4   Column 167   Coefficient 0.00000000
         when "001110100111" => A <= "000000000000000000"; -- Line 4   Column 168   Coefficient 0.00000000
         when "001110101000" => A <= "000000000000000000"; -- Line 4   Column 169   Coefficient 0.00000000
         when "001110101001" => A <= "000000000000000000"; -- Line 4   Column 170   Coefficient 0.00000000
         when "001110101010" => A <= "000000000000000000"; -- Line 4   Column 171   Coefficient 0.00000000
         when "001110101011" => A <= "000000000000000000"; -- Line 4   Column 172   Coefficient 0.00000000
         when "001110101100" => A <= "000000000000000000"; -- Line 4   Column 173   Coefficient 0.00000000
         when "001110101101" => A <= "000000000000000000"; -- Line 4   Column 174   Coefficient 0.00000000
         when "001110101110" => A <= "000000000000000000"; -- Line 4   Column 175   Coefficient 0.00000000
         when "001110101111" => A <= "000000000000000000"; -- Line 4   Column 176   Coefficient 0.00000000
         when "001110110000" => A <= "000000000000000000"; -- Line 4   Column 177   Coefficient 0.00000000
         when "001110110001" => A <= "000000000000000000"; -- Line 4   Column 178   Coefficient 0.00000000
         when "001110110010" => A <= "000000000000000000"; -- Line 4   Column 179   Coefficient 0.00000000
         when "001110110011" => A <= "000000000000000000"; -- Line 4   Column 180   Coefficient 0.00000000
         when "001110110100" => A <= "000000000000000000"; -- Line 4   Column 181   Coefficient 0.00000000
         when "001110110101" => A <= "000000000000000000"; -- Line 4   Column 182   Coefficient 0.00000000
         when "001110110110" => A <= "000000000000000000"; -- Line 4   Column 183   Coefficient 0.00000000
         when "001110110111" => A <= "000000000000000000"; -- Line 4   Column 184   Coefficient 0.00000000
         when "001110111000" => A <= "000000000000000000"; -- Line 4   Column 185   Coefficient 0.00000000
         when "001110111001" => A <= "000000000000000000"; -- Line 4   Column 186   Coefficient 0.00000000
         when "001110111010" => A <= "000000000000000000"; -- Line 4   Column 187   Coefficient 0.00000000
         when "001110111011" => A <= "000000000000000000"; -- Line 4   Column 188   Coefficient 0.00000000
         when "001110111100" => A <= "000000000000000000"; -- Line 4   Column 189   Coefficient 0.00000000
         when "001110111101" => A <= "000000000000000000"; -- Line 4   Column 190   Coefficient 0.00000000
         when "001110111110" => A <= "000000000000000000"; -- Line 4   Column 191   Coefficient 0.00000000
         when "001110111111" => A <= "000000000000000000"; -- Line 4   Column 192   Coefficient 0.00000000
         when "001111000000" => A <= "000000000000000000"; -- Line 4   Column 193   Coefficient 0.00000000
         when "001111000001" => A <= "000000000000000000"; -- Line 4   Column 194   Coefficient 0.00000000
         when "001111000010" => A <= "000000000000000000"; -- Line 4   Column 195   Coefficient 0.00000000
         when "001111000011" => A <= "000000000000000000"; -- Line 4   Column 196   Coefficient 0.00000000
         when "001111000100" => A <= "000000000000000000"; -- Line 4   Column 197   Coefficient 0.00000000
         when "001111000101" => A <= "000000000000000000"; -- Line 4   Column 198   Coefficient 0.00000000
         when "001111000110" => A <= "000000000000000000"; -- Line 4   Column 199   Coefficient 0.00000000
         when "001111000111" => A <= "000000000000000000"; -- Line 4   Column 200   Coefficient 0.00000000
         when "001111001000" => A <= "000000000000000000"; -- Line 4   Column 201   Coefficient 0.00000000
         when "001111001001" => A <= "000000000000000000"; -- Line 4   Column 202   Coefficient 0.00000000
         when "001111001010" => A <= "000000000000000000"; -- Line 4   Column 203   Coefficient 0.00000000
         when "001111001011" => A <= "000000000000000000"; -- Line 4   Column 204   Coefficient 0.00000000
         when "001111001100" => A <= "000000000000000000"; -- Line 4   Column 205   Coefficient 0.00000000
         when "001111001101" => A <= "000000000000000000"; -- Line 4   Column 206   Coefficient 0.00000000
         when "001111001110" => A <= "000000000000000000"; -- Line 4   Column 207   Coefficient 0.00000000
         when "001111001111" => A <= "000000000000000000"; -- Line 4   Column 208   Coefficient 0.00000000
         when "001111010000" => A <= "000000000000000000"; -- Line 4   Column 209   Coefficient 0.00000000
         when "001111010001" => A <= "000000000000000000"; -- Line 4   Column 210   Coefficient 0.00000000
         when "001111010010" => A <= "000000000000000000"; -- Line 4   Column 211   Coefficient 0.00000000
         when "001111010011" => A <= "000000000000000000"; -- Line 4   Column 212   Coefficient 0.00000000
         when "001111010100" => A <= "000000000000000000"; -- Line 4   Column 213   Coefficient 0.00000000
         when "001111010101" => A <= "000000000000000000"; -- Line 4   Column 214   Coefficient 0.00000000
         when "001111010110" => A <= "000000000000000000"; -- Line 4   Column 215   Coefficient 0.00000000
         when "001111010111" => A <= "000000000000000000"; -- Line 4   Column 216   Coefficient 0.00000000
         when "001111011000" => A <= "000000000000000000"; -- Line 4   Column 217   Coefficient 0.00000000
         when "001111011001" => A <= "000000000000000000"; -- Line 4   Column 218   Coefficient 0.00000000
         when "001111011010" => A <= "000000000000000000"; -- Line 4   Column 219   Coefficient 0.00000000
         when "001111011011" => A <= "000000000000000000"; -- Line 4   Column 220   Coefficient 0.00000000
         when "001111011100" => A <= "000000000000000000"; -- Line 4   Column 221   Coefficient 0.00000000
         when "001111011101" => A <= "000000000000000000"; -- Line 4   Column 222   Coefficient 0.00000000
         when "001111011110" => A <= "000000000000000000"; -- Line 4   Column 223   Coefficient 0.00000000
         when "001111011111" => A <= "000000000000000000"; -- Line 4   Column 224   Coefficient 0.00000000
         when "001111100000" => A <= "000000000000000000"; -- Line 4   Column 225   Coefficient 0.00000000
         when "001111100001" => A <= "000000000000000000"; -- Line 4   Column 226   Coefficient 0.00000000
         when "001111100010" => A <= "000000000000000000"; -- Line 4   Column 227   Coefficient 0.00000000
         when "001111100011" => A <= "000000000000000000"; -- Line 4   Column 228   Coefficient 0.00000000
         when "001111100100" => A <= "000000000000000000"; -- Line 4   Column 229   Coefficient 0.00000000
         when "001111100101" => A <= "000000000000000000"; -- Line 4   Column 230   Coefficient 0.00000000
         when "001111100110" => A <= "000000000000000000"; -- Line 4   Column 231   Coefficient 0.00000000
         when "001111100111" => A <= "000000000000000000"; -- Line 4   Column 232   Coefficient 0.00000000
         when "001111101000" => A <= "000000000000000000"; -- Line 4   Column 233   Coefficient 0.00000000
         when "001111101001" => A <= "000000000000000000"; -- Line 4   Column 234   Coefficient 0.00000000
         when "001111101010" => A <= "000000000000000000"; -- Line 4   Column 235   Coefficient 0.00000000
         when "001111101011" => A <= "000000000000000000"; -- Line 4   Column 236   Coefficient 0.00000000
         when "001111101100" => A <= "000000000000000000"; -- Line 4   Column 237   Coefficient 0.00000000
         when "001111101101" => A <= "000000000000000000"; -- Line 4   Column 238   Coefficient 0.00000000
         when "001111101110" => A <= "000000000000000000"; -- Line 4   Column 239   Coefficient 0.00000000
         when "001111101111" => A <= "000000000000000000"; -- Line 4   Column 240   Coefficient 0.00000000
         when "001111110000" => A <= "000000000000000000"; -- Line 4   Column 241   Coefficient 0.00000000
         when "001111110001" => A <= "000000000000000000"; -- Line 4   Column 242   Coefficient 0.00000000
         when "001111110010" => A <= "000000000000000000"; -- Line 4   Column 243   Coefficient 0.00000000
         when "001111110011" => A <= "000000000000000000"; -- Line 4   Column 244   Coefficient 0.00000000
         when "001111110100" => A <= "000000000000000000"; -- Line 4   Column 245   Coefficient 0.00000000
         when "001111110101" => A <= "000000000000000000"; -- Line 4   Column 246   Coefficient 0.00000000
         when "001111110110" => A <= "000000000000000000"; -- Line 4   Column 247   Coefficient 0.00000000
         when "001111110111" => A <= "000000000000000000"; -- Line 4   Column 248   Coefficient 0.00000000
         when "001111111000" => A <= "000000000000000000"; -- Line 4   Column 249   Coefficient 0.00000000
         when "001111111001" => A <= "000000000000000000"; -- Line 4   Column 250   Coefficient 0.00000000
         when "001111111010" => A <= "000000000000000000"; -- Line 4   Column 251   Coefficient 0.00000000
         when "001111111011" => A <= "000000000000000000"; -- Line 4   Column 252   Coefficient 0.00000000
         when "001111111100" => A <= "000000000000000000"; -- Line 4   Column 253   Coefficient 0.00000000
         when "001111111101" => A <= "000000000000000000"; -- Line 4   Column 254   Coefficient 0.00000000
         when "001111111110" => A <= "000000000000000000"; -- Line 4   Column 255   Coefficient 0.00000000
         when "001111111111" => A <= "000000000000000000"; -- Line 4   Column 256   Coefficient 0.00000000
         when "010000000000" => A <= "000000000000000000"; -- Line 5   Column 1   Coefficient 0.00000000
         when "010000000001" => A <= "000000000000000000"; -- Line 5   Column 2   Coefficient 0.00000000
         when "010000000010" => A <= "000000000000000000"; -- Line 5   Column 3   Coefficient 0.00000000
         when "010000000011" => A <= "000000000000000000"; -- Line 5   Column 4   Coefficient 0.00000000
         when "010000000100" => A <= "000000000000000000"; -- Line 5   Column 5   Coefficient 0.00000000
         when "010000000101" => A <= "000000000000000000"; -- Line 5   Column 6   Coefficient 0.00000000
         when "010000000110" => A <= "000000000000000000"; -- Line 5   Column 7   Coefficient 0.00000000
         when "010000000111" => A <= "000000000000000000"; -- Line 5   Column 8   Coefficient 0.00000000
         when "010000001000" => A <= "000000000000000000"; -- Line 5   Column 9   Coefficient 0.00000000
         when "010000001001" => A <= "000000000000000000"; -- Line 5   Column 10   Coefficient 0.00000000
         when "010000001010" => A <= "000000000000000000"; -- Line 5   Column 11   Coefficient 0.00000000
         when "010000001011" => A <= "000000000000000000"; -- Line 5   Column 12   Coefficient 0.00000000
         when "010000001100" => A <= "000000000000000000"; -- Line 5   Column 13   Coefficient 0.00000000
         when "010000001101" => A <= "000000000000000000"; -- Line 5   Column 14   Coefficient 0.00000000
         when "010000001110" => A <= "000000000000000000"; -- Line 5   Column 15   Coefficient 0.00000000
         when "010000001111" => A <= "000000000000000000"; -- Line 5   Column 16   Coefficient 0.00000000
         when "010000010000" => A <= "000000000000000000"; -- Line 5   Column 17   Coefficient 0.00000000
         when "010000010001" => A <= "000000000000000000"; -- Line 5   Column 18   Coefficient 0.00000000
         when "010000010010" => A <= "000000000000000000"; -- Line 5   Column 19   Coefficient 0.00000000
         when "010000010011" => A <= "000000000000000000"; -- Line 5   Column 20   Coefficient 0.00000000
         when "010000010100" => A <= "000000000000000000"; -- Line 5   Column 21   Coefficient 0.00000000
         when "010000010101" => A <= "000000000000000000"; -- Line 5   Column 22   Coefficient 0.00000000
         when "010000010110" => A <= "000000000000000000"; -- Line 5   Column 23   Coefficient 0.00000000
         when "010000010111" => A <= "000000000000000000"; -- Line 5   Column 24   Coefficient 0.00000000
         when "010000011000" => A <= "000000000000000000"; -- Line 5   Column 25   Coefficient 0.00000000
         when "010000011001" => A <= "000000000000000000"; -- Line 5   Column 26   Coefficient 0.00000000
         when "010000011010" => A <= "000000000000000000"; -- Line 5   Column 27   Coefficient 0.00000000
         when "010000011011" => A <= "000000000000000000"; -- Line 5   Column 28   Coefficient 0.00000000
         when "010000011100" => A <= "000000000000000000"; -- Line 5   Column 29   Coefficient 0.00000000
         when "010000011101" => A <= "000000000000000000"; -- Line 5   Column 30   Coefficient 0.00000000
         when "010000011110" => A <= "000000000000000000"; -- Line 5   Column 31   Coefficient 0.00000000
         when "010000011111" => A <= "000000000000000000"; -- Line 5   Column 32   Coefficient 0.00000000
         when "010000100000" => A <= "000000000000000000"; -- Line 5   Column 33   Coefficient 0.00000000
         when "010000100001" => A <= "000000000000000000"; -- Line 5   Column 34   Coefficient 0.00000000
         when "010000100010" => A <= "000000000000000000"; -- Line 5   Column 35   Coefficient 0.00000000
         when "010000100011" => A <= "000000000000000000"; -- Line 5   Column 36   Coefficient 0.00000000
         when "010000100100" => A <= "000000000000000000"; -- Line 5   Column 37   Coefficient 0.00000000
         when "010000100101" => A <= "000000000000000000"; -- Line 5   Column 38   Coefficient 0.00000000
         when "010000100110" => A <= "000000000000000000"; -- Line 5   Column 39   Coefficient 0.00000000
         when "010000100111" => A <= "000000000000000000"; -- Line 5   Column 40   Coefficient 0.00000000
         when "010000101000" => A <= "000000000000000000"; -- Line 5   Column 41   Coefficient 0.00000000
         when "010000101001" => A <= "000000000000000000"; -- Line 5   Column 42   Coefficient 0.00000000
         when "010000101010" => A <= "000000000000000000"; -- Line 5   Column 43   Coefficient 0.00000000
         when "010000101011" => A <= "000000000000000000"; -- Line 5   Column 44   Coefficient 0.00000000
         when "010000101100" => A <= "000000000000000000"; -- Line 5   Column 45   Coefficient 0.00000000
         when "010000101101" => A <= "000000000000000000"; -- Line 5   Column 46   Coefficient 0.00000000
         when "010000101110" => A <= "000000000000000000"; -- Line 5   Column 47   Coefficient 0.00000000
         when "010000101111" => A <= "000000000000000000"; -- Line 5   Column 48   Coefficient 0.00000000
         when "010000110000" => A <= "000000000000000000"; -- Line 5   Column 49   Coefficient 0.00000000
         when "010000110001" => A <= "000000000000000000"; -- Line 5   Column 50   Coefficient 0.00000000
         when "010000110010" => A <= "000000000000000000"; -- Line 5   Column 51   Coefficient 0.00000000
         when "010000110011" => A <= "000000000000000000"; -- Line 5   Column 52   Coefficient 0.00000000
         when "010000110100" => A <= "000000000000000000"; -- Line 5   Column 53   Coefficient 0.00000000
         when "010000110101" => A <= "000000000000000000"; -- Line 5   Column 54   Coefficient 0.00000000
         when "010000110110" => A <= "000000000000000000"; -- Line 5   Column 55   Coefficient 0.00000000
         when "010000110111" => A <= "000000000000000000"; -- Line 5   Column 56   Coefficient 0.00000000
         when "010000111000" => A <= "000000000000000000"; -- Line 5   Column 57   Coefficient 0.00000000
         when "010000111001" => A <= "000000000000000000"; -- Line 5   Column 58   Coefficient 0.00000000
         when "010000111010" => A <= "000000000000000000"; -- Line 5   Column 59   Coefficient 0.00000000
         when "010000111011" => A <= "000000000000000000"; -- Line 5   Column 60   Coefficient 0.00000000
         when "010000111100" => A <= "000000000000000000"; -- Line 5   Column 61   Coefficient 0.00000000
         when "010000111101" => A <= "000000000000000000"; -- Line 5   Column 62   Coefficient 0.00000000
         when "010000111110" => A <= "000000000000000000"; -- Line 5   Column 63   Coefficient 0.00000000
         when "010000111111" => A <= "000000000000000000"; -- Line 5   Column 64   Coefficient 0.00000000
         when "010001000000" => A <= "000000000000001001"; -- Line 5   Column 65   Coefficient 0.00003433
         when "010001000001" => A <= "000000000000000011"; -- Line 5   Column 66   Coefficient 0.00001144
         when "010001000010" => A <= "111111111111001011"; -- Line 5   Column 67   Coefficient -0.00020218
         when "010001000011" => A <= "111111111110100110"; -- Line 5   Column 68   Coefficient -0.00034332
         when "010001000100" => A <= "111111111110010010"; -- Line 5   Column 69   Coefficient -0.00041962
         when "010001000101" => A <= "111111111111010011"; -- Line 5   Column 70   Coefficient -0.00017166
         when "010001000110" => A <= "000000000011111000"; -- Line 5   Column 71   Coefficient 0.00094604
         when "010001000111" => A <= "000000001000010011"; -- Line 5   Column 72   Coefficient 0.00202560
         when "010001001000" => A <= "000000001010110110"; -- Line 5   Column 73   Coefficient 0.00264740
         when "010001001001" => A <= "000000001101001100"; -- Line 5   Column 74   Coefficient 0.00321960
         when "010001001010" => A <= "000000001111111100"; -- Line 5   Column 75   Coefficient 0.00389099
         when "010001001011" => A <= "000000010000011000"; -- Line 5   Column 76   Coefficient 0.00399780
         when "010001001100" => A <= "000000001111000010"; -- Line 5   Column 77   Coefficient 0.00366974
         when "010001001101" => A <= "000000000111011010"; -- Line 5   Column 78   Coefficient 0.00180817
         when "010001001110" => A <= "111111110001010101"; -- Line 5   Column 79   Coefficient -0.00358200
         when "010001001111" => A <= "111111011001111001"; -- Line 5   Column 80   Coefficient -0.00930405
         when "010001010000" => A <= "111111000100111001"; -- Line 5   Column 81   Coefficient -0.01443100
         when "010001010001" => A <= "111110110001100001"; -- Line 5   Column 82   Coefficient -0.01916122
         when "010001010010" => A <= "111110100110010011"; -- Line 5   Column 83   Coefficient -0.02190018
         when "010001010011" => A <= "111110011011111010"; -- Line 5   Column 84   Coefficient -0.02443695
         when "010001010100" => A <= "111110010000110000"; -- Line 5   Column 85   Coefficient -0.02716064
         when "010001010101" => A <= "111110000101010011"; -- Line 5   Column 86   Coefficient -0.02995682
         when "010001010110" => A <= "111101110100001010"; -- Line 5   Column 87   Coefficient -0.03414154
         when "010001010111" => A <= "111101100110110000"; -- Line 5   Column 88   Coefficient -0.03741455
         when "010001011000" => A <= "111101100010101111"; -- Line 5   Column 89   Coefficient -0.03839493
         when "010001011001" => A <= "111101100010001110"; -- Line 5   Column 90   Coefficient -0.03852081
         when "010001011010" => A <= "111101100000101101"; -- Line 5   Column 91   Coefficient -0.03889084
         when "010001011011" => A <= "111101101011101110"; -- Line 5   Column 92   Coefficient -0.03620148
         when "010001011100" => A <= "111110000010011110"; -- Line 5   Column 93   Coefficient -0.03064728
         when "010001011101" => A <= "111110110101100100"; -- Line 5   Column 94   Coefficient -0.01817322
         when "010001011110" => A <= "000000100101011001"; -- Line 5   Column 95   Coefficient 0.00912857
         when "010001011111" => A <= "000010011110111100"; -- Line 5   Column 96   Coefficient 0.03880310
         when "010001100000" => A <= "000100010010000101"; -- Line 5   Column 97   Coefficient 0.06691360
         when "010001100001" => A <= "000110000101110011"; -- Line 5   Column 98   Coefficient 0.09516525
         when "010001100010" => A <= "000111100110110001"; -- Line 5   Column 99   Coefficient 0.11883926
         when "010001100011" => A <= "001001000110101001"; -- Line 5   Column 100   Coefficient 0.14224625
         when "010001100100" => A <= "001010101100000111"; -- Line 5   Column 101   Coefficient 0.16701889
         when "010001100101" => A <= "001100001011101000"; -- Line 5   Column 102   Coefficient 0.19033813
         when "010001100110" => A <= "001101100011111111"; -- Line 5   Column 103   Coefficient 0.21191025
         when "010001100111" => A <= "001110110101010100"; -- Line 5   Column 104   Coefficient 0.23176575
         when "010001101000" => A <= "001111111010100001"; -- Line 5   Column 105   Coefficient 0.24866104
         when "010001101001" => A <= "010000111010100101"; -- Line 5   Column 106   Coefficient 0.26430130
         when "010001101010" => A <= "010010000001100011"; -- Line 5   Column 107   Coefficient 0.28162766
         when "010001101011" => A <= "010010110100110100"; -- Line 5   Column 108   Coefficient 0.29414368
         when "010001101100" => A <= "010011010010100110"; -- Line 5   Column 109   Coefficient 0.30141449
         when "010001101101" => A <= "010011000101100111"; -- Line 5   Column 110   Coefficient 0.29824448
         when "010001101110" => A <= "010001011110001011"; -- Line 5   Column 111   Coefficient 0.27299118
         when "010001101111" => A <= "001111100101110011"; -- Line 5   Column 112   Coefficient 0.24360275
         when "010001110000" => A <= "001101110100101001"; -- Line 5   Column 113   Coefficient 0.21597672
         when "010001110001" => A <= "001011111101111010"; -- Line 5   Column 114   Coefficient 0.18698883
         when "010001110010" => A <= "001010011001111000"; -- Line 5   Column 115   Coefficient 0.16256714
         when "010001110011" => A <= "001000110101000000"; -- Line 5   Column 116   Coefficient 0.13793945
         when "010001110100" => A <= "000111000101010101"; -- Line 5   Column 117   Coefficient 0.11067581
         when "010001110101" => A <= "000101100000010101"; -- Line 5   Column 118   Coefficient 0.08601761
         when "010001110110" => A <= "000100010011001101"; -- Line 5   Column 119   Coefficient 0.06718826
         when "010001110111" => A <= "000011001010010011"; -- Line 5   Column 120   Coefficient 0.04938889
         when "010001111000" => A <= "000010000100001011"; -- Line 5   Column 121   Coefficient 0.03226852
         when "010001111001" => A <= "000000111110100110"; -- Line 5   Column 122   Coefficient 0.01528168
         when "010001111010" => A <= "111111101010001000"; -- Line 5   Column 123   Coefficient -0.00534058
         when "010001111011" => A <= "111110100000101100"; -- Line 5   Column 124   Coefficient -0.02326965
         when "010001111100" => A <= "111101100111001110"; -- Line 5   Column 125   Coefficient -0.03730011
         when "010001111101" => A <= "111101000110110001"; -- Line 5   Column 126   Coefficient -0.04522324
         when "010001111110" => A <= "111101011101101101"; -- Line 5   Column 127   Coefficient -0.03962326
         when "010001111111" => A <= "111101111110110001"; -- Line 5   Column 128   Coefficient -0.03155136
         when "010010000000" => A <= "111110011010010101"; -- Line 5   Column 129   Coefficient -0.02482224
         when "010010000001" => A <= "111110111010000001"; -- Line 5   Column 130   Coefficient -0.01708603
         when "010010000010" => A <= "111111010000101110"; -- Line 5   Column 131   Coefficient -0.01154327
         when "010010000011" => A <= "111111100111100010"; -- Line 5   Column 132   Coefficient -0.00597382
         when "010010000100" => A <= "000000000100100100"; -- Line 5   Column 133   Coefficient 0.00111389
         when "010010000101" => A <= "000000011000110111"; -- Line 5   Column 134   Coefficient 0.00606918
         when "010010000110" => A <= "000000010111101010"; -- Line 5   Column 135   Coefficient 0.00577545
         when "010010000111" => A <= "000000010100111001"; -- Line 5   Column 136   Coefficient 0.00510025
         when "010010001000" => A <= "000000010100110111"; -- Line 5   Column 137   Coefficient 0.00509262
         when "010010001001" => A <= "000000010110010000"; -- Line 5   Column 138   Coefficient 0.00543213
         when "010010001010" => A <= "000000100010100100"; -- Line 5   Column 139   Coefficient 0.00843811
         when "010010001011" => A <= "000000101101010111"; -- Line 5   Column 140   Coefficient 0.01107407
         when "010010001100" => A <= "000000110010101110"; -- Line 5   Column 141   Coefficient 0.01238251
         when "010010001101" => A <= "000000110100010110"; -- Line 5   Column 142   Coefficient 0.01277924
         when "010010001110" => A <= "000000101011110101"; -- Line 5   Column 143   Coefficient 0.01070023
         when "010010001111" => A <= "000000100001110011"; -- Line 5   Column 144   Coefficient 0.00825119
         when "010010010000" => A <= "000000011001110100"; -- Line 5   Column 145   Coefficient 0.00630188
         when "010010010001" => A <= "000000010001001000"; -- Line 5   Column 146   Coefficient 0.00418091
         when "010010010010" => A <= "000000001001011000"; -- Line 5   Column 147   Coefficient 0.00228882
         when "010010010011" => A <= "000000000010010011"; -- Line 5   Column 148   Coefficient 0.00056076
         when "010010010100" => A <= "111111111010111001"; -- Line 5   Column 149   Coefficient -0.00124741
         when "010010010101" => A <= "111111110110011111"; -- Line 5   Column 150   Coefficient -0.00232315
         when "010010010110" => A <= "111111111001000110"; -- Line 5   Column 151   Coefficient -0.00168610
         when "010010010111" => A <= "111111111100011110"; -- Line 5   Column 152   Coefficient -0.00086212
         when "010010011000" => A <= "111111111110110111"; -- Line 5   Column 153   Coefficient -0.00027847
         when "010010011001" => A <= "000000000001001011"; -- Line 5   Column 154   Coefficient 0.00028610
         when "010010011010" => A <= "000000000001001000"; -- Line 5   Column 155   Coefficient 0.00027466
         when "010010011011" => A <= "000000000001000010"; -- Line 5   Column 156   Coefficient 0.00025177
         when "010010011100" => A <= "000000000001111110"; -- Line 5   Column 157   Coefficient 0.00048065
         when "010010011101" => A <= "000000000010010101"; -- Line 5   Column 158   Coefficient 0.00056839
         when "010010011110" => A <= "000000000001100101"; -- Line 5   Column 159   Coefficient 0.00038528
         when "010010011111" => A <= "000000000000110011"; -- Line 5   Column 160   Coefficient 0.00019455
         when "010010100000" => A <= "000000000000000111"; -- Line 5   Column 161   Coefficient 0.00002670
         when "010010100001" => A <= "111111111111100110"; -- Line 5   Column 162   Coefficient -0.00009918
         when "010010100010" => A <= "111111111111110100"; -- Line 5   Column 163   Coefficient -0.00004578
         when "010010100011" => A <= "000000000000000011"; -- Line 5   Column 164   Coefficient 0.00001144
         when "010010100100" => A <= "000000000000000100"; -- Line 5   Column 165   Coefficient 0.00001526
         when "010010100101" => A <= "000000000000000110"; -- Line 5   Column 166   Coefficient 0.00002289
         when "010010100110" => A <= "000000000000000011"; -- Line 5   Column 167   Coefficient 0.00001144
         when "010010100111" => A <= "111111111111111111"; -- Line 5   Column 168   Coefficient -0.00000381
         when "010010101000" => A <= "000000000000000000"; -- Line 5   Column 169   Coefficient 0.00000000
         when "010010101001" => A <= "000000000000000000"; -- Line 5   Column 170   Coefficient 0.00000000
         when "010010101010" => A <= "000000000000000000"; -- Line 5   Column 171   Coefficient 0.00000000
         when "010010101011" => A <= "000000000000000000"; -- Line 5   Column 172   Coefficient 0.00000000
         when "010010101100" => A <= "000000000000000000"; -- Line 5   Column 173   Coefficient 0.00000000
         when "010010101101" => A <= "000000000000000000"; -- Line 5   Column 174   Coefficient 0.00000000
         when "010010101110" => A <= "000000000000000000"; -- Line 5   Column 175   Coefficient 0.00000000
         when "010010101111" => A <= "000000000000000000"; -- Line 5   Column 176   Coefficient 0.00000000
         when "010010110000" => A <= "000000000000000000"; -- Line 5   Column 177   Coefficient 0.00000000
         when "010010110001" => A <= "000000000000000000"; -- Line 5   Column 178   Coefficient 0.00000000
         when "010010110010" => A <= "000000000000000000"; -- Line 5   Column 179   Coefficient 0.00000000
         when "010010110011" => A <= "000000000000000000"; -- Line 5   Column 180   Coefficient 0.00000000
         when "010010110100" => A <= "000000000000000000"; -- Line 5   Column 181   Coefficient 0.00000000
         when "010010110101" => A <= "000000000000000000"; -- Line 5   Column 182   Coefficient 0.00000000
         when "010010110110" => A <= "000000000000000000"; -- Line 5   Column 183   Coefficient 0.00000000
         when "010010110111" => A <= "000000000000000000"; -- Line 5   Column 184   Coefficient 0.00000000
         when "010010111000" => A <= "000000000000000000"; -- Line 5   Column 185   Coefficient 0.00000000
         when "010010111001" => A <= "000000000000000000"; -- Line 5   Column 186   Coefficient 0.00000000
         when "010010111010" => A <= "000000000000000000"; -- Line 5   Column 187   Coefficient 0.00000000
         when "010010111011" => A <= "000000000000000000"; -- Line 5   Column 188   Coefficient 0.00000000
         when "010010111100" => A <= "000000000000000000"; -- Line 5   Column 189   Coefficient 0.00000000
         when "010010111101" => A <= "000000000000000000"; -- Line 5   Column 190   Coefficient 0.00000000
         when "010010111110" => A <= "000000000000000000"; -- Line 5   Column 191   Coefficient 0.00000000
         when "010010111111" => A <= "000000000000000000"; -- Line 5   Column 192   Coefficient 0.00000000
         when "010011000000" => A <= "000000000000000000"; -- Line 5   Column 193   Coefficient 0.00000000
         when "010011000001" => A <= "000000000000000000"; -- Line 5   Column 194   Coefficient 0.00000000
         when "010011000010" => A <= "000000000000000000"; -- Line 5   Column 195   Coefficient 0.00000000
         when "010011000011" => A <= "000000000000000000"; -- Line 5   Column 196   Coefficient 0.00000000
         when "010011000100" => A <= "000000000000000000"; -- Line 5   Column 197   Coefficient 0.00000000
         when "010011000101" => A <= "000000000000000000"; -- Line 5   Column 198   Coefficient 0.00000000
         when "010011000110" => A <= "000000000000000000"; -- Line 5   Column 199   Coefficient 0.00000000
         when "010011000111" => A <= "000000000000000000"; -- Line 5   Column 200   Coefficient 0.00000000
         when "010011001000" => A <= "000000000000000000"; -- Line 5   Column 201   Coefficient 0.00000000
         when "010011001001" => A <= "000000000000000000"; -- Line 5   Column 202   Coefficient 0.00000000
         when "010011001010" => A <= "000000000000000000"; -- Line 5   Column 203   Coefficient 0.00000000
         when "010011001011" => A <= "000000000000000000"; -- Line 5   Column 204   Coefficient 0.00000000
         when "010011001100" => A <= "000000000000000000"; -- Line 5   Column 205   Coefficient 0.00000000
         when "010011001101" => A <= "000000000000000000"; -- Line 5   Column 206   Coefficient 0.00000000
         when "010011001110" => A <= "000000000000000000"; -- Line 5   Column 207   Coefficient 0.00000000
         when "010011001111" => A <= "000000000000000000"; -- Line 5   Column 208   Coefficient 0.00000000
         when "010011010000" => A <= "000000000000000000"; -- Line 5   Column 209   Coefficient 0.00000000
         when "010011010001" => A <= "000000000000000000"; -- Line 5   Column 210   Coefficient 0.00000000
         when "010011010010" => A <= "000000000000000000"; -- Line 5   Column 211   Coefficient 0.00000000
         when "010011010011" => A <= "000000000000000000"; -- Line 5   Column 212   Coefficient 0.00000000
         when "010011010100" => A <= "000000000000000000"; -- Line 5   Column 213   Coefficient 0.00000000
         when "010011010101" => A <= "000000000000000000"; -- Line 5   Column 214   Coefficient 0.00000000
         when "010011010110" => A <= "000000000000000000"; -- Line 5   Column 215   Coefficient 0.00000000
         when "010011010111" => A <= "000000000000000000"; -- Line 5   Column 216   Coefficient 0.00000000
         when "010011011000" => A <= "000000000000000000"; -- Line 5   Column 217   Coefficient 0.00000000
         when "010011011001" => A <= "000000000000000000"; -- Line 5   Column 218   Coefficient 0.00000000
         when "010011011010" => A <= "000000000000000000"; -- Line 5   Column 219   Coefficient 0.00000000
         when "010011011011" => A <= "000000000000000000"; -- Line 5   Column 220   Coefficient 0.00000000
         when "010011011100" => A <= "000000000000000000"; -- Line 5   Column 221   Coefficient 0.00000000
         when "010011011101" => A <= "000000000000000000"; -- Line 5   Column 222   Coefficient 0.00000000
         when "010011011110" => A <= "000000000000000000"; -- Line 5   Column 223   Coefficient 0.00000000
         when "010011011111" => A <= "000000000000000000"; -- Line 5   Column 224   Coefficient 0.00000000
         when "010011100000" => A <= "000000000000000000"; -- Line 5   Column 225   Coefficient 0.00000000
         when "010011100001" => A <= "000000000000000000"; -- Line 5   Column 226   Coefficient 0.00000000
         when "010011100010" => A <= "000000000000000000"; -- Line 5   Column 227   Coefficient 0.00000000
         when "010011100011" => A <= "000000000000000000"; -- Line 5   Column 228   Coefficient 0.00000000
         when "010011100100" => A <= "000000000000000000"; -- Line 5   Column 229   Coefficient 0.00000000
         when "010011100101" => A <= "000000000000000000"; -- Line 5   Column 230   Coefficient 0.00000000
         when "010011100110" => A <= "000000000000000000"; -- Line 5   Column 231   Coefficient 0.00000000
         when "010011100111" => A <= "000000000000000000"; -- Line 5   Column 232   Coefficient 0.00000000
         when "010011101000" => A <= "000000000000000000"; -- Line 5   Column 233   Coefficient 0.00000000
         when "010011101001" => A <= "000000000000000000"; -- Line 5   Column 234   Coefficient 0.00000000
         when "010011101010" => A <= "000000000000000000"; -- Line 5   Column 235   Coefficient 0.00000000
         when "010011101011" => A <= "000000000000000000"; -- Line 5   Column 236   Coefficient 0.00000000
         when "010011101100" => A <= "000000000000000000"; -- Line 5   Column 237   Coefficient 0.00000000
         when "010011101101" => A <= "000000000000000000"; -- Line 5   Column 238   Coefficient 0.00000000
         when "010011101110" => A <= "000000000000000000"; -- Line 5   Column 239   Coefficient 0.00000000
         when "010011101111" => A <= "000000000000000000"; -- Line 5   Column 240   Coefficient 0.00000000
         when "010011110000" => A <= "000000000000000000"; -- Line 5   Column 241   Coefficient 0.00000000
         when "010011110001" => A <= "000000000000000000"; -- Line 5   Column 242   Coefficient 0.00000000
         when "010011110010" => A <= "000000000000000000"; -- Line 5   Column 243   Coefficient 0.00000000
         when "010011110011" => A <= "000000000000000000"; -- Line 5   Column 244   Coefficient 0.00000000
         when "010011110100" => A <= "000000000000000000"; -- Line 5   Column 245   Coefficient 0.00000000
         when "010011110101" => A <= "000000000000000000"; -- Line 5   Column 246   Coefficient 0.00000000
         when "010011110110" => A <= "000000000000000000"; -- Line 5   Column 247   Coefficient 0.00000000
         when "010011110111" => A <= "000000000000000000"; -- Line 5   Column 248   Coefficient 0.00000000
         when "010011111000" => A <= "000000000000000000"; -- Line 5   Column 249   Coefficient 0.00000000
         when "010011111001" => A <= "000000000000000000"; -- Line 5   Column 250   Coefficient 0.00000000
         when "010011111010" => A <= "000000000000000000"; -- Line 5   Column 251   Coefficient 0.00000000
         when "010011111011" => A <= "000000000000000000"; -- Line 5   Column 252   Coefficient 0.00000000
         when "010011111100" => A <= "000000000000000000"; -- Line 5   Column 253   Coefficient 0.00000000
         when "010011111101" => A <= "000000000000000000"; -- Line 5   Column 254   Coefficient 0.00000000
         when "010011111110" => A <= "000000000000000000"; -- Line 5   Column 255   Coefficient 0.00000000
         when "010011111111" => A <= "000000000000000000"; -- Line 5   Column 256   Coefficient 0.00000000
         when "010100000000" => A <= "000000000000000000"; -- Line 6   Column 1   Coefficient 0.00000000
         when "010100000001" => A <= "000000000000000000"; -- Line 6   Column 2   Coefficient 0.00000000
         when "010100000010" => A <= "000000000000000000"; -- Line 6   Column 3   Coefficient 0.00000000
         when "010100000011" => A <= "000000000000000000"; -- Line 6   Column 4   Coefficient 0.00000000
         when "010100000100" => A <= "000000000000000000"; -- Line 6   Column 5   Coefficient 0.00000000
         when "010100000101" => A <= "000000000000000000"; -- Line 6   Column 6   Coefficient 0.00000000
         when "010100000110" => A <= "000000000000000000"; -- Line 6   Column 7   Coefficient 0.00000000
         when "010100000111" => A <= "000000000000000000"; -- Line 6   Column 8   Coefficient 0.00000000
         when "010100001000" => A <= "000000000000000000"; -- Line 6   Column 9   Coefficient 0.00000000
         when "010100001001" => A <= "000000000000000000"; -- Line 6   Column 10   Coefficient 0.00000000
         when "010100001010" => A <= "000000000000000000"; -- Line 6   Column 11   Coefficient 0.00000000
         when "010100001011" => A <= "000000000000000000"; -- Line 6   Column 12   Coefficient 0.00000000
         when "010100001100" => A <= "000000000000000000"; -- Line 6   Column 13   Coefficient 0.00000000
         when "010100001101" => A <= "000000000000000000"; -- Line 6   Column 14   Coefficient 0.00000000
         when "010100001110" => A <= "000000000000000000"; -- Line 6   Column 15   Coefficient 0.00000000
         when "010100001111" => A <= "000000000000000000"; -- Line 6   Column 16   Coefficient 0.00000000
         when "010100010000" => A <= "000000000000000000"; -- Line 6   Column 17   Coefficient 0.00000000
         when "010100010001" => A <= "000000000000000000"; -- Line 6   Column 18   Coefficient 0.00000000
         when "010100010010" => A <= "000000000000000000"; -- Line 6   Column 19   Coefficient 0.00000000
         when "010100010011" => A <= "000000000000000000"; -- Line 6   Column 20   Coefficient 0.00000000
         when "010100010100" => A <= "000000000000000000"; -- Line 6   Column 21   Coefficient 0.00000000
         when "010100010101" => A <= "000000000000000000"; -- Line 6   Column 22   Coefficient 0.00000000
         when "010100010110" => A <= "000000000000000000"; -- Line 6   Column 23   Coefficient 0.00000000
         when "010100010111" => A <= "000000000000000000"; -- Line 6   Column 24   Coefficient 0.00000000
         when "010100011000" => A <= "000000000000000000"; -- Line 6   Column 25   Coefficient 0.00000000
         when "010100011001" => A <= "000000000000000000"; -- Line 6   Column 26   Coefficient 0.00000000
         when "010100011010" => A <= "000000000000000000"; -- Line 6   Column 27   Coefficient 0.00000000
         when "010100011011" => A <= "000000000000000000"; -- Line 6   Column 28   Coefficient 0.00000000
         when "010100011100" => A <= "000000000000000000"; -- Line 6   Column 29   Coefficient 0.00000000
         when "010100011101" => A <= "000000000000000000"; -- Line 6   Column 30   Coefficient 0.00000000
         when "010100011110" => A <= "000000000000000000"; -- Line 6   Column 31   Coefficient 0.00000000
         when "010100011111" => A <= "000000000000000000"; -- Line 6   Column 32   Coefficient 0.00000000
         when "010100100000" => A <= "000000000000000000"; -- Line 6   Column 33   Coefficient 0.00000000
         when "010100100001" => A <= "000000000000000000"; -- Line 6   Column 34   Coefficient 0.00000000
         when "010100100010" => A <= "000000000000000000"; -- Line 6   Column 35   Coefficient 0.00000000
         when "010100100011" => A <= "000000000000000000"; -- Line 6   Column 36   Coefficient 0.00000000
         when "010100100100" => A <= "000000000000000000"; -- Line 6   Column 37   Coefficient 0.00000000
         when "010100100101" => A <= "000000000000000000"; -- Line 6   Column 38   Coefficient 0.00000000
         when "010100100110" => A <= "000000000000000000"; -- Line 6   Column 39   Coefficient 0.00000000
         when "010100100111" => A <= "000000000000000000"; -- Line 6   Column 40   Coefficient 0.00000000
         when "010100101000" => A <= "000000000000000000"; -- Line 6   Column 41   Coefficient 0.00000000
         when "010100101001" => A <= "000000000000000000"; -- Line 6   Column 42   Coefficient 0.00000000
         when "010100101010" => A <= "000000000000000000"; -- Line 6   Column 43   Coefficient 0.00000000
         when "010100101011" => A <= "000000000000000000"; -- Line 6   Column 44   Coefficient 0.00000000
         when "010100101100" => A <= "000000000000000000"; -- Line 6   Column 45   Coefficient 0.00000000
         when "010100101101" => A <= "000000000000000000"; -- Line 6   Column 46   Coefficient 0.00000000
         when "010100101110" => A <= "000000000000000000"; -- Line 6   Column 47   Coefficient 0.00000000
         when "010100101111" => A <= "000000000000000000"; -- Line 6   Column 48   Coefficient 0.00000000
         when "010100110000" => A <= "000000000000000000"; -- Line 6   Column 49   Coefficient 0.00000000
         when "010100110001" => A <= "000000000000000000"; -- Line 6   Column 50   Coefficient 0.00000000
         when "010100110010" => A <= "000000000000000000"; -- Line 6   Column 51   Coefficient 0.00000000
         when "010100110011" => A <= "000000000000000000"; -- Line 6   Column 52   Coefficient 0.00000000
         when "010100110100" => A <= "000000000000000000"; -- Line 6   Column 53   Coefficient 0.00000000
         when "010100110101" => A <= "000000000000000000"; -- Line 6   Column 54   Coefficient 0.00000000
         when "010100110110" => A <= "000000000000000000"; -- Line 6   Column 55   Coefficient 0.00000000
         when "010100110111" => A <= "000000000000000000"; -- Line 6   Column 56   Coefficient 0.00000000
         when "010100111000" => A <= "000000000000000000"; -- Line 6   Column 57   Coefficient 0.00000000
         when "010100111001" => A <= "000000000000000000"; -- Line 6   Column 58   Coefficient 0.00000000
         when "010100111010" => A <= "000000000000000000"; -- Line 6   Column 59   Coefficient 0.00000000
         when "010100111011" => A <= "000000000000000000"; -- Line 6   Column 60   Coefficient 0.00000000
         when "010100111100" => A <= "000000000000000000"; -- Line 6   Column 61   Coefficient 0.00000000
         when "010100111101" => A <= "000000000000000000"; -- Line 6   Column 62   Coefficient 0.00000000
         when "010100111110" => A <= "000000000000000000"; -- Line 6   Column 63   Coefficient 0.00000000
         when "010100111111" => A <= "000000000000000000"; -- Line 6   Column 64   Coefficient 0.00000000
         when "010101000000" => A <= "000000000000000000"; -- Line 6   Column 65   Coefficient 0.00000000
         when "010101000001" => A <= "000000000000000000"; -- Line 6   Column 66   Coefficient 0.00000000
         when "010101000010" => A <= "000000000000000000"; -- Line 6   Column 67   Coefficient 0.00000000
         when "010101000011" => A <= "000000000000000000"; -- Line 6   Column 68   Coefficient 0.00000000
         when "010101000100" => A <= "000000000000000000"; -- Line 6   Column 69   Coefficient 0.00000000
         when "010101000101" => A <= "000000000000000000"; -- Line 6   Column 70   Coefficient 0.00000000
         when "010101000110" => A <= "000000000000000000"; -- Line 6   Column 71   Coefficient 0.00000000
         when "010101000111" => A <= "000000000000000000"; -- Line 6   Column 72   Coefficient 0.00000000
         when "010101001000" => A <= "000000000000000000"; -- Line 6   Column 73   Coefficient 0.00000000
         when "010101001001" => A <= "000000000000000000"; -- Line 6   Column 74   Coefficient 0.00000000
         when "010101001010" => A <= "000000000000000000"; -- Line 6   Column 75   Coefficient 0.00000000
         when "010101001011" => A <= "000000000000000000"; -- Line 6   Column 76   Coefficient 0.00000000
         when "010101001100" => A <= "000000000000000000"; -- Line 6   Column 77   Coefficient 0.00000000
         when "010101001101" => A <= "000000000000000000"; -- Line 6   Column 78   Coefficient 0.00000000
         when "010101001110" => A <= "000000000000000000"; -- Line 6   Column 79   Coefficient 0.00000000
         when "010101001111" => A <= "000000000000000000"; -- Line 6   Column 80   Coefficient 0.00000000
         when "010101010000" => A <= "000000000000001001"; -- Line 6   Column 81   Coefficient 0.00003433
         when "010101010001" => A <= "000000000000000011"; -- Line 6   Column 82   Coefficient 0.00001144
         when "010101010010" => A <= "111111111111001011"; -- Line 6   Column 83   Coefficient -0.00020218
         when "010101010011" => A <= "111111111110100110"; -- Line 6   Column 84   Coefficient -0.00034332
         when "010101010100" => A <= "111111111110010010"; -- Line 6   Column 85   Coefficient -0.00041962
         when "010101010101" => A <= "111111111111010011"; -- Line 6   Column 86   Coefficient -0.00017166
         when "010101010110" => A <= "000000000011111000"; -- Line 6   Column 87   Coefficient 0.00094604
         when "010101010111" => A <= "000000001000010011"; -- Line 6   Column 88   Coefficient 0.00202560
         when "010101011000" => A <= "000000001010110110"; -- Line 6   Column 89   Coefficient 0.00264740
         when "010101011001" => A <= "000000001101001100"; -- Line 6   Column 90   Coefficient 0.00321960
         when "010101011010" => A <= "000000001111111100"; -- Line 6   Column 91   Coefficient 0.00389099
         when "010101011011" => A <= "000000010000011000"; -- Line 6   Column 92   Coefficient 0.00399780
         when "010101011100" => A <= "000000001111000010"; -- Line 6   Column 93   Coefficient 0.00366974
         when "010101011101" => A <= "000000000111011010"; -- Line 6   Column 94   Coefficient 0.00180817
         when "010101011110" => A <= "111111110001010101"; -- Line 6   Column 95   Coefficient -0.00358200
         when "010101011111" => A <= "111111011001111001"; -- Line 6   Column 96   Coefficient -0.00930405
         when "010101100000" => A <= "111111000100111001"; -- Line 6   Column 97   Coefficient -0.01443100
         when "010101100001" => A <= "111110110001100001"; -- Line 6   Column 98   Coefficient -0.01916122
         when "010101100010" => A <= "111110100110010011"; -- Line 6   Column 99   Coefficient -0.02190018
         when "010101100011" => A <= "111110011011111010"; -- Line 6   Column 100   Coefficient -0.02443695
         when "010101100100" => A <= "111110010000110000"; -- Line 6   Column 101   Coefficient -0.02716064
         when "010101100101" => A <= "111110000101010011"; -- Line 6   Column 102   Coefficient -0.02995682
         when "010101100110" => A <= "111101110100001010"; -- Line 6   Column 103   Coefficient -0.03414154
         when "010101100111" => A <= "111101100110110000"; -- Line 6   Column 104   Coefficient -0.03741455
         when "010101101000" => A <= "111101100010101111"; -- Line 6   Column 105   Coefficient -0.03839493
         when "010101101001" => A <= "111101100010001110"; -- Line 6   Column 106   Coefficient -0.03852081
         when "010101101010" => A <= "111101100000101101"; -- Line 6   Column 107   Coefficient -0.03889084
         when "010101101011" => A <= "111101101011101110"; -- Line 6   Column 108   Coefficient -0.03620148
         when "010101101100" => A <= "111110000010011110"; -- Line 6   Column 109   Coefficient -0.03064728
         when "010101101101" => A <= "111110110101100100"; -- Line 6   Column 110   Coefficient -0.01817322
         when "010101101110" => A <= "000000100101011001"; -- Line 6   Column 111   Coefficient 0.00912857
         when "010101101111" => A <= "000010011110111100"; -- Line 6   Column 112   Coefficient 0.03880310
         when "010101110000" => A <= "000100010010000101"; -- Line 6   Column 113   Coefficient 0.06691360
         when "010101110001" => A <= "000110000101110011"; -- Line 6   Column 114   Coefficient 0.09516525
         when "010101110010" => A <= "000111100110110001"; -- Line 6   Column 115   Coefficient 0.11883926
         when "010101110011" => A <= "001001000110101001"; -- Line 6   Column 116   Coefficient 0.14224625
         when "010101110100" => A <= "001010101100000111"; -- Line 6   Column 117   Coefficient 0.16701889
         when "010101110101" => A <= "001100001011101000"; -- Line 6   Column 118   Coefficient 0.19033813
         when "010101110110" => A <= "001101100011111111"; -- Line 6   Column 119   Coefficient 0.21191025
         when "010101110111" => A <= "001110110101010100"; -- Line 6   Column 120   Coefficient 0.23176575
         when "010101111000" => A <= "001111111010100001"; -- Line 6   Column 121   Coefficient 0.24866104
         when "010101111001" => A <= "010000111010100101"; -- Line 6   Column 122   Coefficient 0.26430130
         when "010101111010" => A <= "010010000001100011"; -- Line 6   Column 123   Coefficient 0.28162766
         when "010101111011" => A <= "010010110100110100"; -- Line 6   Column 124   Coefficient 0.29414368
         when "010101111100" => A <= "010011010010100110"; -- Line 6   Column 125   Coefficient 0.30141449
         when "010101111101" => A <= "010011000101100111"; -- Line 6   Column 126   Coefficient 0.29824448
         when "010101111110" => A <= "010001011110001011"; -- Line 6   Column 127   Coefficient 0.27299118
         when "010101111111" => A <= "001111100101110011"; -- Line 6   Column 128   Coefficient 0.24360275
         when "010110000000" => A <= "001101110100101001"; -- Line 6   Column 129   Coefficient 0.21597672
         when "010110000001" => A <= "001011111101111010"; -- Line 6   Column 130   Coefficient 0.18698883
         when "010110000010" => A <= "001010011001111000"; -- Line 6   Column 131   Coefficient 0.16256714
         when "010110000011" => A <= "001000110101000000"; -- Line 6   Column 132   Coefficient 0.13793945
         when "010110000100" => A <= "000111000101010101"; -- Line 6   Column 133   Coefficient 0.11067581
         when "010110000101" => A <= "000101100000010101"; -- Line 6   Column 134   Coefficient 0.08601761
         when "010110000110" => A <= "000100010011001101"; -- Line 6   Column 135   Coefficient 0.06718826
         when "010110000111" => A <= "000011001010010011"; -- Line 6   Column 136   Coefficient 0.04938889
         when "010110001000" => A <= "000010000100001011"; -- Line 6   Column 137   Coefficient 0.03226852
         when "010110001001" => A <= "000000111110100110"; -- Line 6   Column 138   Coefficient 0.01528168
         when "010110001010" => A <= "111111101010001000"; -- Line 6   Column 139   Coefficient -0.00534058
         when "010110001011" => A <= "111110100000101100"; -- Line 6   Column 140   Coefficient -0.02326965
         when "010110001100" => A <= "111101100111001110"; -- Line 6   Column 141   Coefficient -0.03730011
         when "010110001101" => A <= "111101000110110001"; -- Line 6   Column 142   Coefficient -0.04522324
         when "010110001110" => A <= "111101011101101101"; -- Line 6   Column 143   Coefficient -0.03962326
         when "010110001111" => A <= "111101111110110001"; -- Line 6   Column 144   Coefficient -0.03155136
         when "010110010000" => A <= "111110011010010101"; -- Line 6   Column 145   Coefficient -0.02482224
         when "010110010001" => A <= "111110111010000001"; -- Line 6   Column 146   Coefficient -0.01708603
         when "010110010010" => A <= "111111010000101110"; -- Line 6   Column 147   Coefficient -0.01154327
         when "010110010011" => A <= "111111100111100010"; -- Line 6   Column 148   Coefficient -0.00597382
         when "010110010100" => A <= "000000000100100100"; -- Line 6   Column 149   Coefficient 0.00111389
         when "010110010101" => A <= "000000011000110111"; -- Line 6   Column 150   Coefficient 0.00606918
         when "010110010110" => A <= "000000010111101010"; -- Line 6   Column 151   Coefficient 0.00577545
         when "010110010111" => A <= "000000010100111001"; -- Line 6   Column 152   Coefficient 0.00510025
         when "010110011000" => A <= "000000010100110111"; -- Line 6   Column 153   Coefficient 0.00509262
         when "010110011001" => A <= "000000010110010000"; -- Line 6   Column 154   Coefficient 0.00543213
         when "010110011010" => A <= "000000100010100100"; -- Line 6   Column 155   Coefficient 0.00843811
         when "010110011011" => A <= "000000101101010111"; -- Line 6   Column 156   Coefficient 0.01107407
         when "010110011100" => A <= "000000110010101110"; -- Line 6   Column 157   Coefficient 0.01238251
         when "010110011101" => A <= "000000110100010110"; -- Line 6   Column 158   Coefficient 0.01277924
         when "010110011110" => A <= "000000101011110101"; -- Line 6   Column 159   Coefficient 0.01070023
         when "010110011111" => A <= "000000100001110011"; -- Line 6   Column 160   Coefficient 0.00825119
         when "010110100000" => A <= "000000011001110100"; -- Line 6   Column 161   Coefficient 0.00630188
         when "010110100001" => A <= "000000010001001000"; -- Line 6   Column 162   Coefficient 0.00418091
         when "010110100010" => A <= "000000001001011000"; -- Line 6   Column 163   Coefficient 0.00228882
         when "010110100011" => A <= "000000000010010011"; -- Line 6   Column 164   Coefficient 0.00056076
         when "010110100100" => A <= "111111111010111001"; -- Line 6   Column 165   Coefficient -0.00124741
         when "010110100101" => A <= "111111110110011111"; -- Line 6   Column 166   Coefficient -0.00232315
         when "010110100110" => A <= "111111111001000110"; -- Line 6   Column 167   Coefficient -0.00168610
         when "010110100111" => A <= "111111111100011110"; -- Line 6   Column 168   Coefficient -0.00086212
         when "010110101000" => A <= "111111111110110111"; -- Line 6   Column 169   Coefficient -0.00027847
         when "010110101001" => A <= "000000000001001011"; -- Line 6   Column 170   Coefficient 0.00028610
         when "010110101010" => A <= "000000000001001000"; -- Line 6   Column 171   Coefficient 0.00027466
         when "010110101011" => A <= "000000000001000010"; -- Line 6   Column 172   Coefficient 0.00025177
         when "010110101100" => A <= "000000000001111110"; -- Line 6   Column 173   Coefficient 0.00048065
         when "010110101101" => A <= "000000000010010101"; -- Line 6   Column 174   Coefficient 0.00056839
         when "010110101110" => A <= "000000000001100101"; -- Line 6   Column 175   Coefficient 0.00038528
         when "010110101111" => A <= "000000000000110011"; -- Line 6   Column 176   Coefficient 0.00019455
         when "010110110000" => A <= "000000000000000111"; -- Line 6   Column 177   Coefficient 0.00002670
         when "010110110001" => A <= "111111111111100110"; -- Line 6   Column 178   Coefficient -0.00009918
         when "010110110010" => A <= "111111111111110100"; -- Line 6   Column 179   Coefficient -0.00004578
         when "010110110011" => A <= "000000000000000011"; -- Line 6   Column 180   Coefficient 0.00001144
         when "010110110100" => A <= "000000000000000100"; -- Line 6   Column 181   Coefficient 0.00001526
         when "010110110101" => A <= "000000000000000110"; -- Line 6   Column 182   Coefficient 0.00002289
         when "010110110110" => A <= "000000000000000011"; -- Line 6   Column 183   Coefficient 0.00001144
         when "010110110111" => A <= "111111111111111111"; -- Line 6   Column 184   Coefficient -0.00000381
         when "010110111000" => A <= "000000000000000000"; -- Line 6   Column 185   Coefficient 0.00000000
         when "010110111001" => A <= "000000000000000000"; -- Line 6   Column 186   Coefficient 0.00000000
         when "010110111010" => A <= "000000000000000000"; -- Line 6   Column 187   Coefficient 0.00000000
         when "010110111011" => A <= "000000000000000000"; -- Line 6   Column 188   Coefficient 0.00000000
         when "010110111100" => A <= "000000000000000000"; -- Line 6   Column 189   Coefficient 0.00000000
         when "010110111101" => A <= "000000000000000000"; -- Line 6   Column 190   Coefficient 0.00000000
         when "010110111110" => A <= "000000000000000000"; -- Line 6   Column 191   Coefficient 0.00000000
         when "010110111111" => A <= "000000000000000000"; -- Line 6   Column 192   Coefficient 0.00000000
         when "010111000000" => A <= "000000000000000000"; -- Line 6   Column 193   Coefficient 0.00000000
         when "010111000001" => A <= "000000000000000000"; -- Line 6   Column 194   Coefficient 0.00000000
         when "010111000010" => A <= "000000000000000000"; -- Line 6   Column 195   Coefficient 0.00000000
         when "010111000011" => A <= "000000000000000000"; -- Line 6   Column 196   Coefficient 0.00000000
         when "010111000100" => A <= "000000000000000000"; -- Line 6   Column 197   Coefficient 0.00000000
         when "010111000101" => A <= "000000000000000000"; -- Line 6   Column 198   Coefficient 0.00000000
         when "010111000110" => A <= "000000000000000000"; -- Line 6   Column 199   Coefficient 0.00000000
         when "010111000111" => A <= "000000000000000000"; -- Line 6   Column 200   Coefficient 0.00000000
         when "010111001000" => A <= "000000000000000000"; -- Line 6   Column 201   Coefficient 0.00000000
         when "010111001001" => A <= "000000000000000000"; -- Line 6   Column 202   Coefficient 0.00000000
         when "010111001010" => A <= "000000000000000000"; -- Line 6   Column 203   Coefficient 0.00000000
         when "010111001011" => A <= "000000000000000000"; -- Line 6   Column 204   Coefficient 0.00000000
         when "010111001100" => A <= "000000000000000000"; -- Line 6   Column 205   Coefficient 0.00000000
         when "010111001101" => A <= "000000000000000000"; -- Line 6   Column 206   Coefficient 0.00000000
         when "010111001110" => A <= "000000000000000000"; -- Line 6   Column 207   Coefficient 0.00000000
         when "010111001111" => A <= "000000000000000000"; -- Line 6   Column 208   Coefficient 0.00000000
         when "010111010000" => A <= "000000000000000000"; -- Line 6   Column 209   Coefficient 0.00000000
         when "010111010001" => A <= "000000000000000000"; -- Line 6   Column 210   Coefficient 0.00000000
         when "010111010010" => A <= "000000000000000000"; -- Line 6   Column 211   Coefficient 0.00000000
         when "010111010011" => A <= "000000000000000000"; -- Line 6   Column 212   Coefficient 0.00000000
         when "010111010100" => A <= "000000000000000000"; -- Line 6   Column 213   Coefficient 0.00000000
         when "010111010101" => A <= "000000000000000000"; -- Line 6   Column 214   Coefficient 0.00000000
         when "010111010110" => A <= "000000000000000000"; -- Line 6   Column 215   Coefficient 0.00000000
         when "010111010111" => A <= "000000000000000000"; -- Line 6   Column 216   Coefficient 0.00000000
         when "010111011000" => A <= "000000000000000000"; -- Line 6   Column 217   Coefficient 0.00000000
         when "010111011001" => A <= "000000000000000000"; -- Line 6   Column 218   Coefficient 0.00000000
         when "010111011010" => A <= "000000000000000000"; -- Line 6   Column 219   Coefficient 0.00000000
         when "010111011011" => A <= "000000000000000000"; -- Line 6   Column 220   Coefficient 0.00000000
         when "010111011100" => A <= "000000000000000000"; -- Line 6   Column 221   Coefficient 0.00000000
         when "010111011101" => A <= "000000000000000000"; -- Line 6   Column 222   Coefficient 0.00000000
         when "010111011110" => A <= "000000000000000000"; -- Line 6   Column 223   Coefficient 0.00000000
         when "010111011111" => A <= "000000000000000000"; -- Line 6   Column 224   Coefficient 0.00000000
         when "010111100000" => A <= "000000000000000000"; -- Line 6   Column 225   Coefficient 0.00000000
         when "010111100001" => A <= "000000000000000000"; -- Line 6   Column 226   Coefficient 0.00000000
         when "010111100010" => A <= "000000000000000000"; -- Line 6   Column 227   Coefficient 0.00000000
         when "010111100011" => A <= "000000000000000000"; -- Line 6   Column 228   Coefficient 0.00000000
         when "010111100100" => A <= "000000000000000000"; -- Line 6   Column 229   Coefficient 0.00000000
         when "010111100101" => A <= "000000000000000000"; -- Line 6   Column 230   Coefficient 0.00000000
         when "010111100110" => A <= "000000000000000000"; -- Line 6   Column 231   Coefficient 0.00000000
         when "010111100111" => A <= "000000000000000000"; -- Line 6   Column 232   Coefficient 0.00000000
         when "010111101000" => A <= "000000000000000000"; -- Line 6   Column 233   Coefficient 0.00000000
         when "010111101001" => A <= "000000000000000000"; -- Line 6   Column 234   Coefficient 0.00000000
         when "010111101010" => A <= "000000000000000000"; -- Line 6   Column 235   Coefficient 0.00000000
         when "010111101011" => A <= "000000000000000000"; -- Line 6   Column 236   Coefficient 0.00000000
         when "010111101100" => A <= "000000000000000000"; -- Line 6   Column 237   Coefficient 0.00000000
         when "010111101101" => A <= "000000000000000000"; -- Line 6   Column 238   Coefficient 0.00000000
         when "010111101110" => A <= "000000000000000000"; -- Line 6   Column 239   Coefficient 0.00000000
         when "010111101111" => A <= "000000000000000000"; -- Line 6   Column 240   Coefficient 0.00000000
         when "010111110000" => A <= "000000000000000000"; -- Line 6   Column 241   Coefficient 0.00000000
         when "010111110001" => A <= "000000000000000000"; -- Line 6   Column 242   Coefficient 0.00000000
         when "010111110010" => A <= "000000000000000000"; -- Line 6   Column 243   Coefficient 0.00000000
         when "010111110011" => A <= "000000000000000000"; -- Line 6   Column 244   Coefficient 0.00000000
         when "010111110100" => A <= "000000000000000000"; -- Line 6   Column 245   Coefficient 0.00000000
         when "010111110101" => A <= "000000000000000000"; -- Line 6   Column 246   Coefficient 0.00000000
         when "010111110110" => A <= "000000000000000000"; -- Line 6   Column 247   Coefficient 0.00000000
         when "010111110111" => A <= "000000000000000000"; -- Line 6   Column 248   Coefficient 0.00000000
         when "010111111000" => A <= "000000000000000000"; -- Line 6   Column 249   Coefficient 0.00000000
         when "010111111001" => A <= "000000000000000000"; -- Line 6   Column 250   Coefficient 0.00000000
         when "010111111010" => A <= "000000000000000000"; -- Line 6   Column 251   Coefficient 0.00000000
         when "010111111011" => A <= "000000000000000000"; -- Line 6   Column 252   Coefficient 0.00000000
         when "010111111100" => A <= "000000000000000000"; -- Line 6   Column 253   Coefficient 0.00000000
         when "010111111101" => A <= "000000000000000000"; -- Line 6   Column 254   Coefficient 0.00000000
         when "010111111110" => A <= "000000000000000000"; -- Line 6   Column 255   Coefficient 0.00000000
         when "010111111111" => A <= "000000000000000000"; -- Line 6   Column 256   Coefficient 0.00000000
         when "011000000000" => A <= "000000000000000000"; -- Line 7   Column 1   Coefficient 0.00000000
         when "011000000001" => A <= "000000000000000000"; -- Line 7   Column 2   Coefficient 0.00000000
         when "011000000010" => A <= "000000000000000000"; -- Line 7   Column 3   Coefficient 0.00000000
         when "011000000011" => A <= "000000000000000000"; -- Line 7   Column 4   Coefficient 0.00000000
         when "011000000100" => A <= "000000000000000000"; -- Line 7   Column 5   Coefficient 0.00000000
         when "011000000101" => A <= "000000000000000000"; -- Line 7   Column 6   Coefficient 0.00000000
         when "011000000110" => A <= "000000000000000000"; -- Line 7   Column 7   Coefficient 0.00000000
         when "011000000111" => A <= "000000000000000000"; -- Line 7   Column 8   Coefficient 0.00000000
         when "011000001000" => A <= "000000000000000000"; -- Line 7   Column 9   Coefficient 0.00000000
         when "011000001001" => A <= "000000000000000000"; -- Line 7   Column 10   Coefficient 0.00000000
         when "011000001010" => A <= "000000000000000000"; -- Line 7   Column 11   Coefficient 0.00000000
         when "011000001011" => A <= "000000000000000000"; -- Line 7   Column 12   Coefficient 0.00000000
         when "011000001100" => A <= "000000000000000000"; -- Line 7   Column 13   Coefficient 0.00000000
         when "011000001101" => A <= "000000000000000000"; -- Line 7   Column 14   Coefficient 0.00000000
         when "011000001110" => A <= "000000000000000000"; -- Line 7   Column 15   Coefficient 0.00000000
         when "011000001111" => A <= "000000000000000000"; -- Line 7   Column 16   Coefficient 0.00000000
         when "011000010000" => A <= "000000000000000000"; -- Line 7   Column 17   Coefficient 0.00000000
         when "011000010001" => A <= "000000000000000000"; -- Line 7   Column 18   Coefficient 0.00000000
         when "011000010010" => A <= "000000000000000000"; -- Line 7   Column 19   Coefficient 0.00000000
         when "011000010011" => A <= "000000000000000000"; -- Line 7   Column 20   Coefficient 0.00000000
         when "011000010100" => A <= "000000000000000000"; -- Line 7   Column 21   Coefficient 0.00000000
         when "011000010101" => A <= "000000000000000000"; -- Line 7   Column 22   Coefficient 0.00000000
         when "011000010110" => A <= "000000000000000000"; -- Line 7   Column 23   Coefficient 0.00000000
         when "011000010111" => A <= "000000000000000000"; -- Line 7   Column 24   Coefficient 0.00000000
         when "011000011000" => A <= "000000000000000000"; -- Line 7   Column 25   Coefficient 0.00000000
         when "011000011001" => A <= "000000000000000000"; -- Line 7   Column 26   Coefficient 0.00000000
         when "011000011010" => A <= "000000000000000000"; -- Line 7   Column 27   Coefficient 0.00000000
         when "011000011011" => A <= "000000000000000000"; -- Line 7   Column 28   Coefficient 0.00000000
         when "011000011100" => A <= "000000000000000000"; -- Line 7   Column 29   Coefficient 0.00000000
         when "011000011101" => A <= "000000000000000000"; -- Line 7   Column 30   Coefficient 0.00000000
         when "011000011110" => A <= "000000000000000000"; -- Line 7   Column 31   Coefficient 0.00000000
         when "011000011111" => A <= "000000000000000000"; -- Line 7   Column 32   Coefficient 0.00000000
         when "011000100000" => A <= "000000000000000000"; -- Line 7   Column 33   Coefficient 0.00000000
         when "011000100001" => A <= "000000000000000000"; -- Line 7   Column 34   Coefficient 0.00000000
         when "011000100010" => A <= "000000000000000000"; -- Line 7   Column 35   Coefficient 0.00000000
         when "011000100011" => A <= "000000000000000000"; -- Line 7   Column 36   Coefficient 0.00000000
         when "011000100100" => A <= "000000000000000000"; -- Line 7   Column 37   Coefficient 0.00000000
         when "011000100101" => A <= "000000000000000000"; -- Line 7   Column 38   Coefficient 0.00000000
         when "011000100110" => A <= "000000000000000000"; -- Line 7   Column 39   Coefficient 0.00000000
         when "011000100111" => A <= "000000000000000000"; -- Line 7   Column 40   Coefficient 0.00000000
         when "011000101000" => A <= "000000000000000000"; -- Line 7   Column 41   Coefficient 0.00000000
         when "011000101001" => A <= "000000000000000000"; -- Line 7   Column 42   Coefficient 0.00000000
         when "011000101010" => A <= "000000000000000000"; -- Line 7   Column 43   Coefficient 0.00000000
         when "011000101011" => A <= "000000000000000000"; -- Line 7   Column 44   Coefficient 0.00000000
         when "011000101100" => A <= "000000000000000000"; -- Line 7   Column 45   Coefficient 0.00000000
         when "011000101101" => A <= "000000000000000000"; -- Line 7   Column 46   Coefficient 0.00000000
         when "011000101110" => A <= "000000000000000000"; -- Line 7   Column 47   Coefficient 0.00000000
         when "011000101111" => A <= "000000000000000000"; -- Line 7   Column 48   Coefficient 0.00000000
         when "011000110000" => A <= "000000000000000000"; -- Line 7   Column 49   Coefficient 0.00000000
         when "011000110001" => A <= "000000000000000000"; -- Line 7   Column 50   Coefficient 0.00000000
         when "011000110010" => A <= "000000000000000000"; -- Line 7   Column 51   Coefficient 0.00000000
         when "011000110011" => A <= "000000000000000000"; -- Line 7   Column 52   Coefficient 0.00000000
         when "011000110100" => A <= "000000000000000000"; -- Line 7   Column 53   Coefficient 0.00000000
         when "011000110101" => A <= "000000000000000000"; -- Line 7   Column 54   Coefficient 0.00000000
         when "011000110110" => A <= "000000000000000000"; -- Line 7   Column 55   Coefficient 0.00000000
         when "011000110111" => A <= "000000000000000000"; -- Line 7   Column 56   Coefficient 0.00000000
         when "011000111000" => A <= "000000000000000000"; -- Line 7   Column 57   Coefficient 0.00000000
         when "011000111001" => A <= "000000000000000000"; -- Line 7   Column 58   Coefficient 0.00000000
         when "011000111010" => A <= "000000000000000000"; -- Line 7   Column 59   Coefficient 0.00000000
         when "011000111011" => A <= "000000000000000000"; -- Line 7   Column 60   Coefficient 0.00000000
         when "011000111100" => A <= "000000000000000000"; -- Line 7   Column 61   Coefficient 0.00000000
         when "011000111101" => A <= "000000000000000000"; -- Line 7   Column 62   Coefficient 0.00000000
         when "011000111110" => A <= "000000000000000000"; -- Line 7   Column 63   Coefficient 0.00000000
         when "011000111111" => A <= "000000000000000000"; -- Line 7   Column 64   Coefficient 0.00000000
         when "011001000000" => A <= "000000000000000000"; -- Line 7   Column 65   Coefficient 0.00000000
         when "011001000001" => A <= "000000000000000000"; -- Line 7   Column 66   Coefficient 0.00000000
         when "011001000010" => A <= "000000000000000000"; -- Line 7   Column 67   Coefficient 0.00000000
         when "011001000011" => A <= "000000000000000000"; -- Line 7   Column 68   Coefficient 0.00000000
         when "011001000100" => A <= "000000000000000000"; -- Line 7   Column 69   Coefficient 0.00000000
         when "011001000101" => A <= "000000000000000000"; -- Line 7   Column 70   Coefficient 0.00000000
         when "011001000110" => A <= "000000000000000000"; -- Line 7   Column 71   Coefficient 0.00000000
         when "011001000111" => A <= "000000000000000000"; -- Line 7   Column 72   Coefficient 0.00000000
         when "011001001000" => A <= "000000000000000000"; -- Line 7   Column 73   Coefficient 0.00000000
         when "011001001001" => A <= "000000000000000000"; -- Line 7   Column 74   Coefficient 0.00000000
         when "011001001010" => A <= "000000000000000000"; -- Line 7   Column 75   Coefficient 0.00000000
         when "011001001011" => A <= "000000000000000000"; -- Line 7   Column 76   Coefficient 0.00000000
         when "011001001100" => A <= "000000000000000000"; -- Line 7   Column 77   Coefficient 0.00000000
         when "011001001101" => A <= "000000000000000000"; -- Line 7   Column 78   Coefficient 0.00000000
         when "011001001110" => A <= "000000000000000000"; -- Line 7   Column 79   Coefficient 0.00000000
         when "011001001111" => A <= "000000000000000000"; -- Line 7   Column 80   Coefficient 0.00000000
         when "011001010000" => A <= "000000000000000000"; -- Line 7   Column 81   Coefficient 0.00000000
         when "011001010001" => A <= "000000000000000000"; -- Line 7   Column 82   Coefficient 0.00000000
         when "011001010010" => A <= "000000000000000000"; -- Line 7   Column 83   Coefficient 0.00000000
         when "011001010011" => A <= "000000000000000000"; -- Line 7   Column 84   Coefficient 0.00000000
         when "011001010100" => A <= "000000000000000000"; -- Line 7   Column 85   Coefficient 0.00000000
         when "011001010101" => A <= "000000000000000000"; -- Line 7   Column 86   Coefficient 0.00000000
         when "011001010110" => A <= "000000000000000000"; -- Line 7   Column 87   Coefficient 0.00000000
         when "011001010111" => A <= "000000000000000000"; -- Line 7   Column 88   Coefficient 0.00000000
         when "011001011000" => A <= "000000000000000000"; -- Line 7   Column 89   Coefficient 0.00000000
         when "011001011001" => A <= "000000000000000000"; -- Line 7   Column 90   Coefficient 0.00000000
         when "011001011010" => A <= "000000000000000000"; -- Line 7   Column 91   Coefficient 0.00000000
         when "011001011011" => A <= "000000000000000000"; -- Line 7   Column 92   Coefficient 0.00000000
         when "011001011100" => A <= "000000000000000000"; -- Line 7   Column 93   Coefficient 0.00000000
         when "011001011101" => A <= "000000000000000000"; -- Line 7   Column 94   Coefficient 0.00000000
         when "011001011110" => A <= "000000000000000000"; -- Line 7   Column 95   Coefficient 0.00000000
         when "011001011111" => A <= "000000000000000000"; -- Line 7   Column 96   Coefficient 0.00000000
         when "011001100000" => A <= "000000000000001001"; -- Line 7   Column 97   Coefficient 0.00003433
         when "011001100001" => A <= "000000000000000011"; -- Line 7   Column 98   Coefficient 0.00001144
         when "011001100010" => A <= "111111111111001011"; -- Line 7   Column 99   Coefficient -0.00020218
         when "011001100011" => A <= "111111111110100110"; -- Line 7   Column 100   Coefficient -0.00034332
         when "011001100100" => A <= "111111111110010010"; -- Line 7   Column 101   Coefficient -0.00041962
         when "011001100101" => A <= "111111111111010011"; -- Line 7   Column 102   Coefficient -0.00017166
         when "011001100110" => A <= "000000000011111000"; -- Line 7   Column 103   Coefficient 0.00094604
         when "011001100111" => A <= "000000001000010011"; -- Line 7   Column 104   Coefficient 0.00202560
         when "011001101000" => A <= "000000001010110110"; -- Line 7   Column 105   Coefficient 0.00264740
         when "011001101001" => A <= "000000001101001100"; -- Line 7   Column 106   Coefficient 0.00321960
         when "011001101010" => A <= "000000001111111100"; -- Line 7   Column 107   Coefficient 0.00389099
         when "011001101011" => A <= "000000010000011000"; -- Line 7   Column 108   Coefficient 0.00399780
         when "011001101100" => A <= "000000001111000010"; -- Line 7   Column 109   Coefficient 0.00366974
         when "011001101101" => A <= "000000000111011010"; -- Line 7   Column 110   Coefficient 0.00180817
         when "011001101110" => A <= "111111110001010101"; -- Line 7   Column 111   Coefficient -0.00358200
         when "011001101111" => A <= "111111011001111001"; -- Line 7   Column 112   Coefficient -0.00930405
         when "011001110000" => A <= "111111000100111001"; -- Line 7   Column 113   Coefficient -0.01443100
         when "011001110001" => A <= "111110110001100001"; -- Line 7   Column 114   Coefficient -0.01916122
         when "011001110010" => A <= "111110100110010011"; -- Line 7   Column 115   Coefficient -0.02190018
         when "011001110011" => A <= "111110011011111010"; -- Line 7   Column 116   Coefficient -0.02443695
         when "011001110100" => A <= "111110010000110000"; -- Line 7   Column 117   Coefficient -0.02716064
         when "011001110101" => A <= "111110000101010011"; -- Line 7   Column 118   Coefficient -0.02995682
         when "011001110110" => A <= "111101110100001010"; -- Line 7   Column 119   Coefficient -0.03414154
         when "011001110111" => A <= "111101100110110000"; -- Line 7   Column 120   Coefficient -0.03741455
         when "011001111000" => A <= "111101100010101111"; -- Line 7   Column 121   Coefficient -0.03839493
         when "011001111001" => A <= "111101100010001110"; -- Line 7   Column 122   Coefficient -0.03852081
         when "011001111010" => A <= "111101100000101101"; -- Line 7   Column 123   Coefficient -0.03889084
         when "011001111011" => A <= "111101101011101110"; -- Line 7   Column 124   Coefficient -0.03620148
         when "011001111100" => A <= "111110000010011110"; -- Line 7   Column 125   Coefficient -0.03064728
         when "011001111101" => A <= "111110110101100100"; -- Line 7   Column 126   Coefficient -0.01817322
         when "011001111110" => A <= "000000100101011001"; -- Line 7   Column 127   Coefficient 0.00912857
         when "011001111111" => A <= "000010011110111100"; -- Line 7   Column 128   Coefficient 0.03880310
         when "011010000000" => A <= "000100010010000101"; -- Line 7   Column 129   Coefficient 0.06691360
         when "011010000001" => A <= "000110000101110011"; -- Line 7   Column 130   Coefficient 0.09516525
         when "011010000010" => A <= "000111100110110001"; -- Line 7   Column 131   Coefficient 0.11883926
         when "011010000011" => A <= "001001000110101001"; -- Line 7   Column 132   Coefficient 0.14224625
         when "011010000100" => A <= "001010101100000111"; -- Line 7   Column 133   Coefficient 0.16701889
         when "011010000101" => A <= "001100001011101000"; -- Line 7   Column 134   Coefficient 0.19033813
         when "011010000110" => A <= "001101100011111111"; -- Line 7   Column 135   Coefficient 0.21191025
         when "011010000111" => A <= "001110110101010100"; -- Line 7   Column 136   Coefficient 0.23176575
         when "011010001000" => A <= "001111111010100001"; -- Line 7   Column 137   Coefficient 0.24866104
         when "011010001001" => A <= "010000111010100101"; -- Line 7   Column 138   Coefficient 0.26430130
         when "011010001010" => A <= "010010000001100011"; -- Line 7   Column 139   Coefficient 0.28162766
         when "011010001011" => A <= "010010110100110100"; -- Line 7   Column 140   Coefficient 0.29414368
         when "011010001100" => A <= "010011010010100110"; -- Line 7   Column 141   Coefficient 0.30141449
         when "011010001101" => A <= "010011000101100111"; -- Line 7   Column 142   Coefficient 0.29824448
         when "011010001110" => A <= "010001011110001011"; -- Line 7   Column 143   Coefficient 0.27299118
         when "011010001111" => A <= "001111100101110011"; -- Line 7   Column 144   Coefficient 0.24360275
         when "011010010000" => A <= "001101110100101001"; -- Line 7   Column 145   Coefficient 0.21597672
         when "011010010001" => A <= "001011111101111010"; -- Line 7   Column 146   Coefficient 0.18698883
         when "011010010010" => A <= "001010011001111000"; -- Line 7   Column 147   Coefficient 0.16256714
         when "011010010011" => A <= "001000110101000000"; -- Line 7   Column 148   Coefficient 0.13793945
         when "011010010100" => A <= "000111000101010101"; -- Line 7   Column 149   Coefficient 0.11067581
         when "011010010101" => A <= "000101100000010101"; -- Line 7   Column 150   Coefficient 0.08601761
         when "011010010110" => A <= "000100010011001101"; -- Line 7   Column 151   Coefficient 0.06718826
         when "011010010111" => A <= "000011001010010011"; -- Line 7   Column 152   Coefficient 0.04938889
         when "011010011000" => A <= "000010000100001011"; -- Line 7   Column 153   Coefficient 0.03226852
         when "011010011001" => A <= "000000111110100110"; -- Line 7   Column 154   Coefficient 0.01528168
         when "011010011010" => A <= "111111101010001000"; -- Line 7   Column 155   Coefficient -0.00534058
         when "011010011011" => A <= "111110100000101100"; -- Line 7   Column 156   Coefficient -0.02326965
         when "011010011100" => A <= "111101100111001110"; -- Line 7   Column 157   Coefficient -0.03730011
         when "011010011101" => A <= "111101000110110001"; -- Line 7   Column 158   Coefficient -0.04522324
         when "011010011110" => A <= "111101011101101101"; -- Line 7   Column 159   Coefficient -0.03962326
         when "011010011111" => A <= "111101111110110001"; -- Line 7   Column 160   Coefficient -0.03155136
         when "011010100000" => A <= "111110011010010101"; -- Line 7   Column 161   Coefficient -0.02482224
         when "011010100001" => A <= "111110111010000001"; -- Line 7   Column 162   Coefficient -0.01708603
         when "011010100010" => A <= "111111010000101110"; -- Line 7   Column 163   Coefficient -0.01154327
         when "011010100011" => A <= "111111100111100010"; -- Line 7   Column 164   Coefficient -0.00597382
         when "011010100100" => A <= "000000000100100100"; -- Line 7   Column 165   Coefficient 0.00111389
         when "011010100101" => A <= "000000011000110111"; -- Line 7   Column 166   Coefficient 0.00606918
         when "011010100110" => A <= "000000010111101010"; -- Line 7   Column 167   Coefficient 0.00577545
         when "011010100111" => A <= "000000010100111001"; -- Line 7   Column 168   Coefficient 0.00510025
         when "011010101000" => A <= "000000010100110111"; -- Line 7   Column 169   Coefficient 0.00509262
         when "011010101001" => A <= "000000010110010000"; -- Line 7   Column 170   Coefficient 0.00543213
         when "011010101010" => A <= "000000100010100100"; -- Line 7   Column 171   Coefficient 0.00843811
         when "011010101011" => A <= "000000101101010111"; -- Line 7   Column 172   Coefficient 0.01107407
         when "011010101100" => A <= "000000110010101110"; -- Line 7   Column 173   Coefficient 0.01238251
         when "011010101101" => A <= "000000110100010110"; -- Line 7   Column 174   Coefficient 0.01277924
         when "011010101110" => A <= "000000101011110101"; -- Line 7   Column 175   Coefficient 0.01070023
         when "011010101111" => A <= "000000100001110011"; -- Line 7   Column 176   Coefficient 0.00825119
         when "011010110000" => A <= "000000011001110100"; -- Line 7   Column 177   Coefficient 0.00630188
         when "011010110001" => A <= "000000010001001000"; -- Line 7   Column 178   Coefficient 0.00418091
         when "011010110010" => A <= "000000001001011000"; -- Line 7   Column 179   Coefficient 0.00228882
         when "011010110011" => A <= "000000000010010011"; -- Line 7   Column 180   Coefficient 0.00056076
         when "011010110100" => A <= "111111111010111001"; -- Line 7   Column 181   Coefficient -0.00124741
         when "011010110101" => A <= "111111110110011111"; -- Line 7   Column 182   Coefficient -0.00232315
         when "011010110110" => A <= "111111111001000110"; -- Line 7   Column 183   Coefficient -0.00168610
         when "011010110111" => A <= "111111111100011110"; -- Line 7   Column 184   Coefficient -0.00086212
         when "011010111000" => A <= "111111111110110111"; -- Line 7   Column 185   Coefficient -0.00027847
         when "011010111001" => A <= "000000000001001011"; -- Line 7   Column 186   Coefficient 0.00028610
         when "011010111010" => A <= "000000000001001000"; -- Line 7   Column 187   Coefficient 0.00027466
         when "011010111011" => A <= "000000000001000010"; -- Line 7   Column 188   Coefficient 0.00025177
         when "011010111100" => A <= "000000000001111110"; -- Line 7   Column 189   Coefficient 0.00048065
         when "011010111101" => A <= "000000000010010101"; -- Line 7   Column 190   Coefficient 0.00056839
         when "011010111110" => A <= "000000000001100101"; -- Line 7   Column 191   Coefficient 0.00038528
         when "011010111111" => A <= "000000000000110011"; -- Line 7   Column 192   Coefficient 0.00019455
         when "011011000000" => A <= "000000000000000111"; -- Line 7   Column 193   Coefficient 0.00002670
         when "011011000001" => A <= "111111111111100110"; -- Line 7   Column 194   Coefficient -0.00009918
         when "011011000010" => A <= "111111111111110100"; -- Line 7   Column 195   Coefficient -0.00004578
         when "011011000011" => A <= "000000000000000011"; -- Line 7   Column 196   Coefficient 0.00001144
         when "011011000100" => A <= "000000000000000100"; -- Line 7   Column 197   Coefficient 0.00001526
         when "011011000101" => A <= "000000000000000110"; -- Line 7   Column 198   Coefficient 0.00002289
         when "011011000110" => A <= "000000000000000011"; -- Line 7   Column 199   Coefficient 0.00001144
         when "011011000111" => A <= "111111111111111111"; -- Line 7   Column 200   Coefficient -0.00000381
         when "011011001000" => A <= "000000000000000000"; -- Line 7   Column 201   Coefficient 0.00000000
         when "011011001001" => A <= "000000000000000000"; -- Line 7   Column 202   Coefficient 0.00000000
         when "011011001010" => A <= "000000000000000000"; -- Line 7   Column 203   Coefficient 0.00000000
         when "011011001011" => A <= "000000000000000000"; -- Line 7   Column 204   Coefficient 0.00000000
         when "011011001100" => A <= "000000000000000000"; -- Line 7   Column 205   Coefficient 0.00000000
         when "011011001101" => A <= "000000000000000000"; -- Line 7   Column 206   Coefficient 0.00000000
         when "011011001110" => A <= "000000000000000000"; -- Line 7   Column 207   Coefficient 0.00000000
         when "011011001111" => A <= "000000000000000000"; -- Line 7   Column 208   Coefficient 0.00000000
         when "011011010000" => A <= "000000000000000000"; -- Line 7   Column 209   Coefficient 0.00000000
         when "011011010001" => A <= "000000000000000000"; -- Line 7   Column 210   Coefficient 0.00000000
         when "011011010010" => A <= "000000000000000000"; -- Line 7   Column 211   Coefficient 0.00000000
         when "011011010011" => A <= "000000000000000000"; -- Line 7   Column 212   Coefficient 0.00000000
         when "011011010100" => A <= "000000000000000000"; -- Line 7   Column 213   Coefficient 0.00000000
         when "011011010101" => A <= "000000000000000000"; -- Line 7   Column 214   Coefficient 0.00000000
         when "011011010110" => A <= "000000000000000000"; -- Line 7   Column 215   Coefficient 0.00000000
         when "011011010111" => A <= "000000000000000000"; -- Line 7   Column 216   Coefficient 0.00000000
         when "011011011000" => A <= "000000000000000000"; -- Line 7   Column 217   Coefficient 0.00000000
         when "011011011001" => A <= "000000000000000000"; -- Line 7   Column 218   Coefficient 0.00000000
         when "011011011010" => A <= "000000000000000000"; -- Line 7   Column 219   Coefficient 0.00000000
         when "011011011011" => A <= "000000000000000000"; -- Line 7   Column 220   Coefficient 0.00000000
         when "011011011100" => A <= "000000000000000000"; -- Line 7   Column 221   Coefficient 0.00000000
         when "011011011101" => A <= "000000000000000000"; -- Line 7   Column 222   Coefficient 0.00000000
         when "011011011110" => A <= "000000000000000000"; -- Line 7   Column 223   Coefficient 0.00000000
         when "011011011111" => A <= "000000000000000000"; -- Line 7   Column 224   Coefficient 0.00000000
         when "011011100000" => A <= "000000000000000000"; -- Line 7   Column 225   Coefficient 0.00000000
         when "011011100001" => A <= "000000000000000000"; -- Line 7   Column 226   Coefficient 0.00000000
         when "011011100010" => A <= "000000000000000000"; -- Line 7   Column 227   Coefficient 0.00000000
         when "011011100011" => A <= "000000000000000000"; -- Line 7   Column 228   Coefficient 0.00000000
         when "011011100100" => A <= "000000000000000000"; -- Line 7   Column 229   Coefficient 0.00000000
         when "011011100101" => A <= "000000000000000000"; -- Line 7   Column 230   Coefficient 0.00000000
         when "011011100110" => A <= "000000000000000000"; -- Line 7   Column 231   Coefficient 0.00000000
         when "011011100111" => A <= "000000000000000000"; -- Line 7   Column 232   Coefficient 0.00000000
         when "011011101000" => A <= "000000000000000000"; -- Line 7   Column 233   Coefficient 0.00000000
         when "011011101001" => A <= "000000000000000000"; -- Line 7   Column 234   Coefficient 0.00000000
         when "011011101010" => A <= "000000000000000000"; -- Line 7   Column 235   Coefficient 0.00000000
         when "011011101011" => A <= "000000000000000000"; -- Line 7   Column 236   Coefficient 0.00000000
         when "011011101100" => A <= "000000000000000000"; -- Line 7   Column 237   Coefficient 0.00000000
         when "011011101101" => A <= "000000000000000000"; -- Line 7   Column 238   Coefficient 0.00000000
         when "011011101110" => A <= "000000000000000000"; -- Line 7   Column 239   Coefficient 0.00000000
         when "011011101111" => A <= "000000000000000000"; -- Line 7   Column 240   Coefficient 0.00000000
         when "011011110000" => A <= "000000000000000000"; -- Line 7   Column 241   Coefficient 0.00000000
         when "011011110001" => A <= "000000000000000000"; -- Line 7   Column 242   Coefficient 0.00000000
         when "011011110010" => A <= "000000000000000000"; -- Line 7   Column 243   Coefficient 0.00000000
         when "011011110011" => A <= "000000000000000000"; -- Line 7   Column 244   Coefficient 0.00000000
         when "011011110100" => A <= "000000000000000000"; -- Line 7   Column 245   Coefficient 0.00000000
         when "011011110101" => A <= "000000000000000000"; -- Line 7   Column 246   Coefficient 0.00000000
         when "011011110110" => A <= "000000000000000000"; -- Line 7   Column 247   Coefficient 0.00000000
         when "011011110111" => A <= "000000000000000000"; -- Line 7   Column 248   Coefficient 0.00000000
         when "011011111000" => A <= "000000000000000000"; -- Line 7   Column 249   Coefficient 0.00000000
         when "011011111001" => A <= "000000000000000000"; -- Line 7   Column 250   Coefficient 0.00000000
         when "011011111010" => A <= "000000000000000000"; -- Line 7   Column 251   Coefficient 0.00000000
         when "011011111011" => A <= "000000000000000000"; -- Line 7   Column 252   Coefficient 0.00000000
         when "011011111100" => A <= "000000000000000000"; -- Line 7   Column 253   Coefficient 0.00000000
         when "011011111101" => A <= "000000000000000000"; -- Line 7   Column 254   Coefficient 0.00000000
         when "011011111110" => A <= "000000000000000000"; -- Line 7   Column 255   Coefficient 0.00000000
         when "011011111111" => A <= "000000000000000000"; -- Line 7   Column 256   Coefficient 0.00000000
         when "011100000000" => A <= "000000000000000000"; -- Line 8   Column 1   Coefficient 0.00000000
         when "011100000001" => A <= "000000000000000000"; -- Line 8   Column 2   Coefficient 0.00000000
         when "011100000010" => A <= "000000000000000000"; -- Line 8   Column 3   Coefficient 0.00000000
         when "011100000011" => A <= "000000000000000000"; -- Line 8   Column 4   Coefficient 0.00000000
         when "011100000100" => A <= "000000000000000000"; -- Line 8   Column 5   Coefficient 0.00000000
         when "011100000101" => A <= "000000000000000000"; -- Line 8   Column 6   Coefficient 0.00000000
         when "011100000110" => A <= "000000000000000000"; -- Line 8   Column 7   Coefficient 0.00000000
         when "011100000111" => A <= "000000000000000000"; -- Line 8   Column 8   Coefficient 0.00000000
         when "011100001000" => A <= "000000000000000000"; -- Line 8   Column 9   Coefficient 0.00000000
         when "011100001001" => A <= "000000000000000000"; -- Line 8   Column 10   Coefficient 0.00000000
         when "011100001010" => A <= "000000000000000000"; -- Line 8   Column 11   Coefficient 0.00000000
         when "011100001011" => A <= "000000000000000000"; -- Line 8   Column 12   Coefficient 0.00000000
         when "011100001100" => A <= "000000000000000000"; -- Line 8   Column 13   Coefficient 0.00000000
         when "011100001101" => A <= "000000000000000000"; -- Line 8   Column 14   Coefficient 0.00000000
         when "011100001110" => A <= "000000000000000000"; -- Line 8   Column 15   Coefficient 0.00000000
         when "011100001111" => A <= "000000000000000000"; -- Line 8   Column 16   Coefficient 0.00000000
         when "011100010000" => A <= "000000000000000000"; -- Line 8   Column 17   Coefficient 0.00000000
         when "011100010001" => A <= "000000000000000000"; -- Line 8   Column 18   Coefficient 0.00000000
         when "011100010010" => A <= "000000000000000000"; -- Line 8   Column 19   Coefficient 0.00000000
         when "011100010011" => A <= "000000000000000000"; -- Line 8   Column 20   Coefficient 0.00000000
         when "011100010100" => A <= "000000000000000000"; -- Line 8   Column 21   Coefficient 0.00000000
         when "011100010101" => A <= "000000000000000000"; -- Line 8   Column 22   Coefficient 0.00000000
         when "011100010110" => A <= "000000000000000000"; -- Line 8   Column 23   Coefficient 0.00000000
         when "011100010111" => A <= "000000000000000000"; -- Line 8   Column 24   Coefficient 0.00000000
         when "011100011000" => A <= "000000000000000000"; -- Line 8   Column 25   Coefficient 0.00000000
         when "011100011001" => A <= "000000000000000000"; -- Line 8   Column 26   Coefficient 0.00000000
         when "011100011010" => A <= "000000000000000000"; -- Line 8   Column 27   Coefficient 0.00000000
         when "011100011011" => A <= "000000000000000000"; -- Line 8   Column 28   Coefficient 0.00000000
         when "011100011100" => A <= "000000000000000000"; -- Line 8   Column 29   Coefficient 0.00000000
         when "011100011101" => A <= "000000000000000000"; -- Line 8   Column 30   Coefficient 0.00000000
         when "011100011110" => A <= "000000000000000000"; -- Line 8   Column 31   Coefficient 0.00000000
         when "011100011111" => A <= "000000000000000000"; -- Line 8   Column 32   Coefficient 0.00000000
         when "011100100000" => A <= "000000000000000000"; -- Line 8   Column 33   Coefficient 0.00000000
         when "011100100001" => A <= "000000000000000000"; -- Line 8   Column 34   Coefficient 0.00000000
         when "011100100010" => A <= "000000000000000000"; -- Line 8   Column 35   Coefficient 0.00000000
         when "011100100011" => A <= "000000000000000000"; -- Line 8   Column 36   Coefficient 0.00000000
         when "011100100100" => A <= "000000000000000000"; -- Line 8   Column 37   Coefficient 0.00000000
         when "011100100101" => A <= "000000000000000000"; -- Line 8   Column 38   Coefficient 0.00000000
         when "011100100110" => A <= "000000000000000000"; -- Line 8   Column 39   Coefficient 0.00000000
         when "011100100111" => A <= "000000000000000000"; -- Line 8   Column 40   Coefficient 0.00000000
         when "011100101000" => A <= "000000000000000000"; -- Line 8   Column 41   Coefficient 0.00000000
         when "011100101001" => A <= "000000000000000000"; -- Line 8   Column 42   Coefficient 0.00000000
         when "011100101010" => A <= "000000000000000000"; -- Line 8   Column 43   Coefficient 0.00000000
         when "011100101011" => A <= "000000000000000000"; -- Line 8   Column 44   Coefficient 0.00000000
         when "011100101100" => A <= "000000000000000000"; -- Line 8   Column 45   Coefficient 0.00000000
         when "011100101101" => A <= "000000000000000000"; -- Line 8   Column 46   Coefficient 0.00000000
         when "011100101110" => A <= "000000000000000000"; -- Line 8   Column 47   Coefficient 0.00000000
         when "011100101111" => A <= "000000000000000000"; -- Line 8   Column 48   Coefficient 0.00000000
         when "011100110000" => A <= "000000000000000000"; -- Line 8   Column 49   Coefficient 0.00000000
         when "011100110001" => A <= "000000000000000000"; -- Line 8   Column 50   Coefficient 0.00000000
         when "011100110010" => A <= "000000000000000000"; -- Line 8   Column 51   Coefficient 0.00000000
         when "011100110011" => A <= "000000000000000000"; -- Line 8   Column 52   Coefficient 0.00000000
         when "011100110100" => A <= "000000000000000000"; -- Line 8   Column 53   Coefficient 0.00000000
         when "011100110101" => A <= "000000000000000000"; -- Line 8   Column 54   Coefficient 0.00000000
         when "011100110110" => A <= "000000000000000000"; -- Line 8   Column 55   Coefficient 0.00000000
         when "011100110111" => A <= "000000000000000000"; -- Line 8   Column 56   Coefficient 0.00000000
         when "011100111000" => A <= "000000000000000000"; -- Line 8   Column 57   Coefficient 0.00000000
         when "011100111001" => A <= "000000000000000000"; -- Line 8   Column 58   Coefficient 0.00000000
         when "011100111010" => A <= "000000000000000000"; -- Line 8   Column 59   Coefficient 0.00000000
         when "011100111011" => A <= "000000000000000000"; -- Line 8   Column 60   Coefficient 0.00000000
         when "011100111100" => A <= "000000000000000000"; -- Line 8   Column 61   Coefficient 0.00000000
         when "011100111101" => A <= "000000000000000000"; -- Line 8   Column 62   Coefficient 0.00000000
         when "011100111110" => A <= "000000000000000000"; -- Line 8   Column 63   Coefficient 0.00000000
         when "011100111111" => A <= "000000000000000000"; -- Line 8   Column 64   Coefficient 0.00000000
         when "011101000000" => A <= "000000000000000000"; -- Line 8   Column 65   Coefficient 0.00000000
         when "011101000001" => A <= "000000000000000000"; -- Line 8   Column 66   Coefficient 0.00000000
         when "011101000010" => A <= "000000000000000000"; -- Line 8   Column 67   Coefficient 0.00000000
         when "011101000011" => A <= "000000000000000000"; -- Line 8   Column 68   Coefficient 0.00000000
         when "011101000100" => A <= "000000000000000000"; -- Line 8   Column 69   Coefficient 0.00000000
         when "011101000101" => A <= "000000000000000000"; -- Line 8   Column 70   Coefficient 0.00000000
         when "011101000110" => A <= "000000000000000000"; -- Line 8   Column 71   Coefficient 0.00000000
         when "011101000111" => A <= "000000000000000000"; -- Line 8   Column 72   Coefficient 0.00000000
         when "011101001000" => A <= "000000000000000000"; -- Line 8   Column 73   Coefficient 0.00000000
         when "011101001001" => A <= "000000000000000000"; -- Line 8   Column 74   Coefficient 0.00000000
         when "011101001010" => A <= "000000000000000000"; -- Line 8   Column 75   Coefficient 0.00000000
         when "011101001011" => A <= "000000000000000000"; -- Line 8   Column 76   Coefficient 0.00000000
         when "011101001100" => A <= "000000000000000000"; -- Line 8   Column 77   Coefficient 0.00000000
         when "011101001101" => A <= "000000000000000000"; -- Line 8   Column 78   Coefficient 0.00000000
         when "011101001110" => A <= "000000000000000000"; -- Line 8   Column 79   Coefficient 0.00000000
         when "011101001111" => A <= "000000000000000000"; -- Line 8   Column 80   Coefficient 0.00000000
         when "011101010000" => A <= "000000000000000000"; -- Line 8   Column 81   Coefficient 0.00000000
         when "011101010001" => A <= "000000000000000000"; -- Line 8   Column 82   Coefficient 0.00000000
         when "011101010010" => A <= "000000000000000000"; -- Line 8   Column 83   Coefficient 0.00000000
         when "011101010011" => A <= "000000000000000000"; -- Line 8   Column 84   Coefficient 0.00000000
         when "011101010100" => A <= "000000000000000000"; -- Line 8   Column 85   Coefficient 0.00000000
         when "011101010101" => A <= "000000000000000000"; -- Line 8   Column 86   Coefficient 0.00000000
         when "011101010110" => A <= "000000000000000000"; -- Line 8   Column 87   Coefficient 0.00000000
         when "011101010111" => A <= "000000000000000000"; -- Line 8   Column 88   Coefficient 0.00000000
         when "011101011000" => A <= "000000000000000000"; -- Line 8   Column 89   Coefficient 0.00000000
         when "011101011001" => A <= "000000000000000000"; -- Line 8   Column 90   Coefficient 0.00000000
         when "011101011010" => A <= "000000000000000000"; -- Line 8   Column 91   Coefficient 0.00000000
         when "011101011011" => A <= "000000000000000000"; -- Line 8   Column 92   Coefficient 0.00000000
         when "011101011100" => A <= "000000000000000000"; -- Line 8   Column 93   Coefficient 0.00000000
         when "011101011101" => A <= "000000000000000000"; -- Line 8   Column 94   Coefficient 0.00000000
         when "011101011110" => A <= "000000000000000000"; -- Line 8   Column 95   Coefficient 0.00000000
         when "011101011111" => A <= "000000000000000000"; -- Line 8   Column 96   Coefficient 0.00000000
         when "011101100000" => A <= "000000000000000000"; -- Line 8   Column 97   Coefficient 0.00000000
         when "011101100001" => A <= "000000000000000000"; -- Line 8   Column 98   Coefficient 0.00000000
         when "011101100010" => A <= "000000000000000000"; -- Line 8   Column 99   Coefficient 0.00000000
         when "011101100011" => A <= "000000000000000000"; -- Line 8   Column 100   Coefficient 0.00000000
         when "011101100100" => A <= "000000000000000000"; -- Line 8   Column 101   Coefficient 0.00000000
         when "011101100101" => A <= "000000000000000000"; -- Line 8   Column 102   Coefficient 0.00000000
         when "011101100110" => A <= "000000000000000000"; -- Line 8   Column 103   Coefficient 0.00000000
         when "011101100111" => A <= "000000000000000000"; -- Line 8   Column 104   Coefficient 0.00000000
         when "011101101000" => A <= "000000000000000000"; -- Line 8   Column 105   Coefficient 0.00000000
         when "011101101001" => A <= "000000000000000000"; -- Line 8   Column 106   Coefficient 0.00000000
         when "011101101010" => A <= "000000000000000000"; -- Line 8   Column 107   Coefficient 0.00000000
         when "011101101011" => A <= "000000000000000000"; -- Line 8   Column 108   Coefficient 0.00000000
         when "011101101100" => A <= "000000000000000000"; -- Line 8   Column 109   Coefficient 0.00000000
         when "011101101101" => A <= "000000000000000000"; -- Line 8   Column 110   Coefficient 0.00000000
         when "011101101110" => A <= "000000000000000000"; -- Line 8   Column 111   Coefficient 0.00000000
         when "011101101111" => A <= "000000000000000000"; -- Line 8   Column 112   Coefficient 0.00000000
         when "011101110000" => A <= "000000000000001001"; -- Line 8   Column 113   Coefficient 0.00003433
         when "011101110001" => A <= "000000000000000011"; -- Line 8   Column 114   Coefficient 0.00001144
         when "011101110010" => A <= "111111111111001011"; -- Line 8   Column 115   Coefficient -0.00020218
         when "011101110011" => A <= "111111111110100110"; -- Line 8   Column 116   Coefficient -0.00034332
         when "011101110100" => A <= "111111111110010010"; -- Line 8   Column 117   Coefficient -0.00041962
         when "011101110101" => A <= "111111111111010011"; -- Line 8   Column 118   Coefficient -0.00017166
         when "011101110110" => A <= "000000000011111000"; -- Line 8   Column 119   Coefficient 0.00094604
         when "011101110111" => A <= "000000001000010011"; -- Line 8   Column 120   Coefficient 0.00202560
         when "011101111000" => A <= "000000001010110110"; -- Line 8   Column 121   Coefficient 0.00264740
         when "011101111001" => A <= "000000001101001100"; -- Line 8   Column 122   Coefficient 0.00321960
         when "011101111010" => A <= "000000001111111100"; -- Line 8   Column 123   Coefficient 0.00389099
         when "011101111011" => A <= "000000010000011000"; -- Line 8   Column 124   Coefficient 0.00399780
         when "011101111100" => A <= "000000001111000010"; -- Line 8   Column 125   Coefficient 0.00366974
         when "011101111101" => A <= "000000000111011010"; -- Line 8   Column 126   Coefficient 0.00180817
         when "011101111110" => A <= "111111110001010101"; -- Line 8   Column 127   Coefficient -0.00358200
         when "011101111111" => A <= "111111011001111001"; -- Line 8   Column 128   Coefficient -0.00930405
         when "011110000000" => A <= "111111000100111001"; -- Line 8   Column 129   Coefficient -0.01443100
         when "011110000001" => A <= "111110110001100001"; -- Line 8   Column 130   Coefficient -0.01916122
         when "011110000010" => A <= "111110100110010011"; -- Line 8   Column 131   Coefficient -0.02190018
         when "011110000011" => A <= "111110011011111010"; -- Line 8   Column 132   Coefficient -0.02443695
         when "011110000100" => A <= "111110010000110000"; -- Line 8   Column 133   Coefficient -0.02716064
         when "011110000101" => A <= "111110000101010011"; -- Line 8   Column 134   Coefficient -0.02995682
         when "011110000110" => A <= "111101110100001010"; -- Line 8   Column 135   Coefficient -0.03414154
         when "011110000111" => A <= "111101100110110000"; -- Line 8   Column 136   Coefficient -0.03741455
         when "011110001000" => A <= "111101100010101111"; -- Line 8   Column 137   Coefficient -0.03839493
         when "011110001001" => A <= "111101100010001110"; -- Line 8   Column 138   Coefficient -0.03852081
         when "011110001010" => A <= "111101100000101101"; -- Line 8   Column 139   Coefficient -0.03889084
         when "011110001011" => A <= "111101101011101110"; -- Line 8   Column 140   Coefficient -0.03620148
         when "011110001100" => A <= "111110000010011110"; -- Line 8   Column 141   Coefficient -0.03064728
         when "011110001101" => A <= "111110110101100100"; -- Line 8   Column 142   Coefficient -0.01817322
         when "011110001110" => A <= "000000100101011001"; -- Line 8   Column 143   Coefficient 0.00912857
         when "011110001111" => A <= "000010011110111100"; -- Line 8   Column 144   Coefficient 0.03880310
         when "011110010000" => A <= "000100010010000101"; -- Line 8   Column 145   Coefficient 0.06691360
         when "011110010001" => A <= "000110000101110011"; -- Line 8   Column 146   Coefficient 0.09516525
         when "011110010010" => A <= "000111100110110001"; -- Line 8   Column 147   Coefficient 0.11883926
         when "011110010011" => A <= "001001000110101001"; -- Line 8   Column 148   Coefficient 0.14224625
         when "011110010100" => A <= "001010101100000111"; -- Line 8   Column 149   Coefficient 0.16701889
         when "011110010101" => A <= "001100001011101000"; -- Line 8   Column 150   Coefficient 0.19033813
         when "011110010110" => A <= "001101100011111111"; -- Line 8   Column 151   Coefficient 0.21191025
         when "011110010111" => A <= "001110110101010100"; -- Line 8   Column 152   Coefficient 0.23176575
         when "011110011000" => A <= "001111111010100001"; -- Line 8   Column 153   Coefficient 0.24866104
         when "011110011001" => A <= "010000111010100101"; -- Line 8   Column 154   Coefficient 0.26430130
         when "011110011010" => A <= "010010000001100011"; -- Line 8   Column 155   Coefficient 0.28162766
         when "011110011011" => A <= "010010110100110100"; -- Line 8   Column 156   Coefficient 0.29414368
         when "011110011100" => A <= "010011010010100110"; -- Line 8   Column 157   Coefficient 0.30141449
         when "011110011101" => A <= "010011000101100111"; -- Line 8   Column 158   Coefficient 0.29824448
         when "011110011110" => A <= "010001011110001011"; -- Line 8   Column 159   Coefficient 0.27299118
         when "011110011111" => A <= "001111100101110011"; -- Line 8   Column 160   Coefficient 0.24360275
         when "011110100000" => A <= "001101110100101001"; -- Line 8   Column 161   Coefficient 0.21597672
         when "011110100001" => A <= "001011111101111010"; -- Line 8   Column 162   Coefficient 0.18698883
         when "011110100010" => A <= "001010011001111000"; -- Line 8   Column 163   Coefficient 0.16256714
         when "011110100011" => A <= "001000110101000000"; -- Line 8   Column 164   Coefficient 0.13793945
         when "011110100100" => A <= "000111000101010101"; -- Line 8   Column 165   Coefficient 0.11067581
         when "011110100101" => A <= "000101100000010101"; -- Line 8   Column 166   Coefficient 0.08601761
         when "011110100110" => A <= "000100010011001101"; -- Line 8   Column 167   Coefficient 0.06718826
         when "011110100111" => A <= "000011001010010011"; -- Line 8   Column 168   Coefficient 0.04938889
         when "011110101000" => A <= "000010000100001011"; -- Line 8   Column 169   Coefficient 0.03226852
         when "011110101001" => A <= "000000111110100110"; -- Line 8   Column 170   Coefficient 0.01528168
         when "011110101010" => A <= "111111101010001000"; -- Line 8   Column 171   Coefficient -0.00534058
         when "011110101011" => A <= "111110100000101100"; -- Line 8   Column 172   Coefficient -0.02326965
         when "011110101100" => A <= "111101100111001110"; -- Line 8   Column 173   Coefficient -0.03730011
         when "011110101101" => A <= "111101000110110001"; -- Line 8   Column 174   Coefficient -0.04522324
         when "011110101110" => A <= "111101011101101101"; -- Line 8   Column 175   Coefficient -0.03962326
         when "011110101111" => A <= "111101111110110001"; -- Line 8   Column 176   Coefficient -0.03155136
         when "011110110000" => A <= "111110011010010101"; -- Line 8   Column 177   Coefficient -0.02482224
         when "011110110001" => A <= "111110111010000001"; -- Line 8   Column 178   Coefficient -0.01708603
         when "011110110010" => A <= "111111010000101110"; -- Line 8   Column 179   Coefficient -0.01154327
         when "011110110011" => A <= "111111100111100010"; -- Line 8   Column 180   Coefficient -0.00597382
         when "011110110100" => A <= "000000000100100100"; -- Line 8   Column 181   Coefficient 0.00111389
         when "011110110101" => A <= "000000011000110111"; -- Line 8   Column 182   Coefficient 0.00606918
         when "011110110110" => A <= "000000010111101010"; -- Line 8   Column 183   Coefficient 0.00577545
         when "011110110111" => A <= "000000010100111001"; -- Line 8   Column 184   Coefficient 0.00510025
         when "011110111000" => A <= "000000010100110111"; -- Line 8   Column 185   Coefficient 0.00509262
         when "011110111001" => A <= "000000010110010000"; -- Line 8   Column 186   Coefficient 0.00543213
         when "011110111010" => A <= "000000100010100100"; -- Line 8   Column 187   Coefficient 0.00843811
         when "011110111011" => A <= "000000101101010111"; -- Line 8   Column 188   Coefficient 0.01107407
         when "011110111100" => A <= "000000110010101110"; -- Line 8   Column 189   Coefficient 0.01238251
         when "011110111101" => A <= "000000110100010110"; -- Line 8   Column 190   Coefficient 0.01277924
         when "011110111110" => A <= "000000101011110101"; -- Line 8   Column 191   Coefficient 0.01070023
         when "011110111111" => A <= "000000100001110011"; -- Line 8   Column 192   Coefficient 0.00825119
         when "011111000000" => A <= "000000011001110100"; -- Line 8   Column 193   Coefficient 0.00630188
         when "011111000001" => A <= "000000010001001000"; -- Line 8   Column 194   Coefficient 0.00418091
         when "011111000010" => A <= "000000001001011000"; -- Line 8   Column 195   Coefficient 0.00228882
         when "011111000011" => A <= "000000000010010011"; -- Line 8   Column 196   Coefficient 0.00056076
         when "011111000100" => A <= "111111111010111001"; -- Line 8   Column 197   Coefficient -0.00124741
         when "011111000101" => A <= "111111110110011111"; -- Line 8   Column 198   Coefficient -0.00232315
         when "011111000110" => A <= "111111111001000110"; -- Line 8   Column 199   Coefficient -0.00168610
         when "011111000111" => A <= "111111111100011110"; -- Line 8   Column 200   Coefficient -0.00086212
         when "011111001000" => A <= "111111111110110111"; -- Line 8   Column 201   Coefficient -0.00027847
         when "011111001001" => A <= "000000000001001011"; -- Line 8   Column 202   Coefficient 0.00028610
         when "011111001010" => A <= "000000000001001000"; -- Line 8   Column 203   Coefficient 0.00027466
         when "011111001011" => A <= "000000000001000010"; -- Line 8   Column 204   Coefficient 0.00025177
         when "011111001100" => A <= "000000000001111110"; -- Line 8   Column 205   Coefficient 0.00048065
         when "011111001101" => A <= "000000000010010101"; -- Line 8   Column 206   Coefficient 0.00056839
         when "011111001110" => A <= "000000000001100101"; -- Line 8   Column 207   Coefficient 0.00038528
         when "011111001111" => A <= "000000000000110011"; -- Line 8   Column 208   Coefficient 0.00019455
         when "011111010000" => A <= "000000000000000111"; -- Line 8   Column 209   Coefficient 0.00002670
         when "011111010001" => A <= "111111111111100110"; -- Line 8   Column 210   Coefficient -0.00009918
         when "011111010010" => A <= "111111111111110100"; -- Line 8   Column 211   Coefficient -0.00004578
         when "011111010011" => A <= "000000000000000011"; -- Line 8   Column 212   Coefficient 0.00001144
         when "011111010100" => A <= "000000000000000100"; -- Line 8   Column 213   Coefficient 0.00001526
         when "011111010101" => A <= "000000000000000110"; -- Line 8   Column 214   Coefficient 0.00002289
         when "011111010110" => A <= "000000000000000011"; -- Line 8   Column 215   Coefficient 0.00001144
         when "011111010111" => A <= "111111111111111111"; -- Line 8   Column 216   Coefficient -0.00000381
         when "011111011000" => A <= "000000000000000000"; -- Line 8   Column 217   Coefficient 0.00000000
         when "011111011001" => A <= "000000000000000000"; -- Line 8   Column 218   Coefficient 0.00000000
         when "011111011010" => A <= "000000000000000000"; -- Line 8   Column 219   Coefficient 0.00000000
         when "011111011011" => A <= "000000000000000000"; -- Line 8   Column 220   Coefficient 0.00000000
         when "011111011100" => A <= "000000000000000000"; -- Line 8   Column 221   Coefficient 0.00000000
         when "011111011101" => A <= "000000000000000000"; -- Line 8   Column 222   Coefficient 0.00000000
         when "011111011110" => A <= "000000000000000000"; -- Line 8   Column 223   Coefficient 0.00000000
         when "011111011111" => A <= "000000000000000000"; -- Line 8   Column 224   Coefficient 0.00000000
         when "011111100000" => A <= "000000000000000000"; -- Line 8   Column 225   Coefficient 0.00000000
         when "011111100001" => A <= "000000000000000000"; -- Line 8   Column 226   Coefficient 0.00000000
         when "011111100010" => A <= "000000000000000000"; -- Line 8   Column 227   Coefficient 0.00000000
         when "011111100011" => A <= "000000000000000000"; -- Line 8   Column 228   Coefficient 0.00000000
         when "011111100100" => A <= "000000000000000000"; -- Line 8   Column 229   Coefficient 0.00000000
         when "011111100101" => A <= "000000000000000000"; -- Line 8   Column 230   Coefficient 0.00000000
         when "011111100110" => A <= "000000000000000000"; -- Line 8   Column 231   Coefficient 0.00000000
         when "011111100111" => A <= "000000000000000000"; -- Line 8   Column 232   Coefficient 0.00000000
         when "011111101000" => A <= "000000000000000000"; -- Line 8   Column 233   Coefficient 0.00000000
         when "011111101001" => A <= "000000000000000000"; -- Line 8   Column 234   Coefficient 0.00000000
         when "011111101010" => A <= "000000000000000000"; -- Line 8   Column 235   Coefficient 0.00000000
         when "011111101011" => A <= "000000000000000000"; -- Line 8   Column 236   Coefficient 0.00000000
         when "011111101100" => A <= "000000000000000000"; -- Line 8   Column 237   Coefficient 0.00000000
         when "011111101101" => A <= "000000000000000000"; -- Line 8   Column 238   Coefficient 0.00000000
         when "011111101110" => A <= "000000000000000000"; -- Line 8   Column 239   Coefficient 0.00000000
         when "011111101111" => A <= "000000000000000000"; -- Line 8   Column 240   Coefficient 0.00000000
         when "011111110000" => A <= "000000000000000000"; -- Line 8   Column 241   Coefficient 0.00000000
         when "011111110001" => A <= "000000000000000000"; -- Line 8   Column 242   Coefficient 0.00000000
         when "011111110010" => A <= "000000000000000000"; -- Line 8   Column 243   Coefficient 0.00000000
         when "011111110011" => A <= "000000000000000000"; -- Line 8   Column 244   Coefficient 0.00000000
         when "011111110100" => A <= "000000000000000000"; -- Line 8   Column 245   Coefficient 0.00000000
         when "011111110101" => A <= "000000000000000000"; -- Line 8   Column 246   Coefficient 0.00000000
         when "011111110110" => A <= "000000000000000000"; -- Line 8   Column 247   Coefficient 0.00000000
         when "011111110111" => A <= "000000000000000000"; -- Line 8   Column 248   Coefficient 0.00000000
         when "011111111000" => A <= "000000000000000000"; -- Line 8   Column 249   Coefficient 0.00000000
         when "011111111001" => A <= "000000000000000000"; -- Line 8   Column 250   Coefficient 0.00000000
         when "011111111010" => A <= "000000000000000000"; -- Line 8   Column 251   Coefficient 0.00000000
         when "011111111011" => A <= "000000000000000000"; -- Line 8   Column 252   Coefficient 0.00000000
         when "011111111100" => A <= "000000000000000000"; -- Line 8   Column 253   Coefficient 0.00000000
         when "011111111101" => A <= "000000000000000000"; -- Line 8   Column 254   Coefficient 0.00000000
         when "011111111110" => A <= "000000000000000000"; -- Line 8   Column 255   Coefficient 0.00000000
         when "011111111111" => A <= "000000000000000000"; -- Line 8   Column 256   Coefficient 0.00000000
         when "100000000000" => A <= "000000000000000000"; -- Line 9   Column 1   Coefficient 0.00000000
         when "100000000001" => A <= "000000000000000000"; -- Line 9   Column 2   Coefficient 0.00000000
         when "100000000010" => A <= "000000000000000000"; -- Line 9   Column 3   Coefficient 0.00000000
         when "100000000011" => A <= "000000000000000000"; -- Line 9   Column 4   Coefficient 0.00000000
         when "100000000100" => A <= "000000000000000000"; -- Line 9   Column 5   Coefficient 0.00000000
         when "100000000101" => A <= "000000000000000000"; -- Line 9   Column 6   Coefficient 0.00000000
         when "100000000110" => A <= "000000000000000000"; -- Line 9   Column 7   Coefficient 0.00000000
         when "100000000111" => A <= "000000000000000000"; -- Line 9   Column 8   Coefficient 0.00000000
         when "100000001000" => A <= "000000000000000000"; -- Line 9   Column 9   Coefficient 0.00000000
         when "100000001001" => A <= "000000000000000000"; -- Line 9   Column 10   Coefficient 0.00000000
         when "100000001010" => A <= "000000000000000000"; -- Line 9   Column 11   Coefficient 0.00000000
         when "100000001011" => A <= "000000000000000000"; -- Line 9   Column 12   Coefficient 0.00000000
         when "100000001100" => A <= "000000000000000000"; -- Line 9   Column 13   Coefficient 0.00000000
         when "100000001101" => A <= "000000000000000000"; -- Line 9   Column 14   Coefficient 0.00000000
         when "100000001110" => A <= "000000000000000000"; -- Line 9   Column 15   Coefficient 0.00000000
         when "100000001111" => A <= "000000000000000000"; -- Line 9   Column 16   Coefficient 0.00000000
         when "100000010000" => A <= "000000000000000000"; -- Line 9   Column 17   Coefficient 0.00000000
         when "100000010001" => A <= "000000000000000000"; -- Line 9   Column 18   Coefficient 0.00000000
         when "100000010010" => A <= "000000000000000000"; -- Line 9   Column 19   Coefficient 0.00000000
         when "100000010011" => A <= "000000000000000000"; -- Line 9   Column 20   Coefficient 0.00000000
         when "100000010100" => A <= "000000000000000000"; -- Line 9   Column 21   Coefficient 0.00000000
         when "100000010101" => A <= "000000000000000000"; -- Line 9   Column 22   Coefficient 0.00000000
         when "100000010110" => A <= "000000000000000000"; -- Line 9   Column 23   Coefficient 0.00000000
         when "100000010111" => A <= "000000000000000000"; -- Line 9   Column 24   Coefficient 0.00000000
         when "100000011000" => A <= "000000000000000000"; -- Line 9   Column 25   Coefficient 0.00000000
         when "100000011001" => A <= "000000000000000000"; -- Line 9   Column 26   Coefficient 0.00000000
         when "100000011010" => A <= "000000000000000000"; -- Line 9   Column 27   Coefficient 0.00000000
         when "100000011011" => A <= "000000000000000000"; -- Line 9   Column 28   Coefficient 0.00000000
         when "100000011100" => A <= "000000000000000000"; -- Line 9   Column 29   Coefficient 0.00000000
         when "100000011101" => A <= "000000000000000000"; -- Line 9   Column 30   Coefficient 0.00000000
         when "100000011110" => A <= "000000000000000000"; -- Line 9   Column 31   Coefficient 0.00000000
         when "100000011111" => A <= "000000000000000000"; -- Line 9   Column 32   Coefficient 0.00000000
         when "100000100000" => A <= "000000000000000000"; -- Line 9   Column 33   Coefficient 0.00000000
         when "100000100001" => A <= "000000000000000000"; -- Line 9   Column 34   Coefficient 0.00000000
         when "100000100010" => A <= "000000000000000000"; -- Line 9   Column 35   Coefficient 0.00000000
         when "100000100011" => A <= "000000000000000000"; -- Line 9   Column 36   Coefficient 0.00000000
         when "100000100100" => A <= "000000000000000000"; -- Line 9   Column 37   Coefficient 0.00000000
         when "100000100101" => A <= "000000000000000000"; -- Line 9   Column 38   Coefficient 0.00000000
         when "100000100110" => A <= "000000000000000000"; -- Line 9   Column 39   Coefficient 0.00000000
         when "100000100111" => A <= "000000000000000000"; -- Line 9   Column 40   Coefficient 0.00000000
         when "100000101000" => A <= "000000000000000000"; -- Line 9   Column 41   Coefficient 0.00000000
         when "100000101001" => A <= "000000000000000000"; -- Line 9   Column 42   Coefficient 0.00000000
         when "100000101010" => A <= "000000000000000000"; -- Line 9   Column 43   Coefficient 0.00000000
         when "100000101011" => A <= "000000000000000000"; -- Line 9   Column 44   Coefficient 0.00000000
         when "100000101100" => A <= "000000000000000000"; -- Line 9   Column 45   Coefficient 0.00000000
         when "100000101101" => A <= "000000000000000000"; -- Line 9   Column 46   Coefficient 0.00000000
         when "100000101110" => A <= "000000000000000000"; -- Line 9   Column 47   Coefficient 0.00000000
         when "100000101111" => A <= "000000000000000000"; -- Line 9   Column 48   Coefficient 0.00000000
         when "100000110000" => A <= "000000000000000000"; -- Line 9   Column 49   Coefficient 0.00000000
         when "100000110001" => A <= "000000000000000000"; -- Line 9   Column 50   Coefficient 0.00000000
         when "100000110010" => A <= "000000000000000000"; -- Line 9   Column 51   Coefficient 0.00000000
         when "100000110011" => A <= "000000000000000000"; -- Line 9   Column 52   Coefficient 0.00000000
         when "100000110100" => A <= "000000000000000000"; -- Line 9   Column 53   Coefficient 0.00000000
         when "100000110101" => A <= "000000000000000000"; -- Line 9   Column 54   Coefficient 0.00000000
         when "100000110110" => A <= "000000000000000000"; -- Line 9   Column 55   Coefficient 0.00000000
         when "100000110111" => A <= "000000000000000000"; -- Line 9   Column 56   Coefficient 0.00000000
         when "100000111000" => A <= "000000000000000000"; -- Line 9   Column 57   Coefficient 0.00000000
         when "100000111001" => A <= "000000000000000000"; -- Line 9   Column 58   Coefficient 0.00000000
         when "100000111010" => A <= "000000000000000000"; -- Line 9   Column 59   Coefficient 0.00000000
         when "100000111011" => A <= "000000000000000000"; -- Line 9   Column 60   Coefficient 0.00000000
         when "100000111100" => A <= "000000000000000000"; -- Line 9   Column 61   Coefficient 0.00000000
         when "100000111101" => A <= "000000000000000000"; -- Line 9   Column 62   Coefficient 0.00000000
         when "100000111110" => A <= "000000000000000000"; -- Line 9   Column 63   Coefficient 0.00000000
         when "100000111111" => A <= "000000000000000000"; -- Line 9   Column 64   Coefficient 0.00000000
         when "100001000000" => A <= "000000000000000000"; -- Line 9   Column 65   Coefficient 0.00000000
         when "100001000001" => A <= "000000000000000000"; -- Line 9   Column 66   Coefficient 0.00000000
         when "100001000010" => A <= "000000000000000000"; -- Line 9   Column 67   Coefficient 0.00000000
         when "100001000011" => A <= "000000000000000000"; -- Line 9   Column 68   Coefficient 0.00000000
         when "100001000100" => A <= "000000000000000000"; -- Line 9   Column 69   Coefficient 0.00000000
         when "100001000101" => A <= "000000000000000000"; -- Line 9   Column 70   Coefficient 0.00000000
         when "100001000110" => A <= "000000000000000000"; -- Line 9   Column 71   Coefficient 0.00000000
         when "100001000111" => A <= "000000000000000000"; -- Line 9   Column 72   Coefficient 0.00000000
         when "100001001000" => A <= "000000000000000000"; -- Line 9   Column 73   Coefficient 0.00000000
         when "100001001001" => A <= "000000000000000000"; -- Line 9   Column 74   Coefficient 0.00000000
         when "100001001010" => A <= "000000000000000000"; -- Line 9   Column 75   Coefficient 0.00000000
         when "100001001011" => A <= "000000000000000000"; -- Line 9   Column 76   Coefficient 0.00000000
         when "100001001100" => A <= "000000000000000000"; -- Line 9   Column 77   Coefficient 0.00000000
         when "100001001101" => A <= "000000000000000000"; -- Line 9   Column 78   Coefficient 0.00000000
         when "100001001110" => A <= "000000000000000000"; -- Line 9   Column 79   Coefficient 0.00000000
         when "100001001111" => A <= "000000000000000000"; -- Line 9   Column 80   Coefficient 0.00000000
         when "100001010000" => A <= "000000000000000000"; -- Line 9   Column 81   Coefficient 0.00000000
         when "100001010001" => A <= "000000000000000000"; -- Line 9   Column 82   Coefficient 0.00000000
         when "100001010010" => A <= "000000000000000000"; -- Line 9   Column 83   Coefficient 0.00000000
         when "100001010011" => A <= "000000000000000000"; -- Line 9   Column 84   Coefficient 0.00000000
         when "100001010100" => A <= "000000000000000000"; -- Line 9   Column 85   Coefficient 0.00000000
         when "100001010101" => A <= "000000000000000000"; -- Line 9   Column 86   Coefficient 0.00000000
         when "100001010110" => A <= "000000000000000000"; -- Line 9   Column 87   Coefficient 0.00000000
         when "100001010111" => A <= "000000000000000000"; -- Line 9   Column 88   Coefficient 0.00000000
         when "100001011000" => A <= "000000000000000000"; -- Line 9   Column 89   Coefficient 0.00000000
         when "100001011001" => A <= "000000000000000000"; -- Line 9   Column 90   Coefficient 0.00000000
         when "100001011010" => A <= "000000000000000000"; -- Line 9   Column 91   Coefficient 0.00000000
         when "100001011011" => A <= "000000000000000000"; -- Line 9   Column 92   Coefficient 0.00000000
         when "100001011100" => A <= "000000000000000000"; -- Line 9   Column 93   Coefficient 0.00000000
         when "100001011101" => A <= "000000000000000000"; -- Line 9   Column 94   Coefficient 0.00000000
         when "100001011110" => A <= "000000000000000000"; -- Line 9   Column 95   Coefficient 0.00000000
         when "100001011111" => A <= "000000000000000000"; -- Line 9   Column 96   Coefficient 0.00000000
         when "100001100000" => A <= "000000000000000000"; -- Line 9   Column 97   Coefficient 0.00000000
         when "100001100001" => A <= "000000000000000000"; -- Line 9   Column 98   Coefficient 0.00000000
         when "100001100010" => A <= "000000000000000000"; -- Line 9   Column 99   Coefficient 0.00000000
         when "100001100011" => A <= "000000000000000000"; -- Line 9   Column 100   Coefficient 0.00000000
         when "100001100100" => A <= "000000000000000000"; -- Line 9   Column 101   Coefficient 0.00000000
         when "100001100101" => A <= "000000000000000000"; -- Line 9   Column 102   Coefficient 0.00000000
         when "100001100110" => A <= "000000000000000000"; -- Line 9   Column 103   Coefficient 0.00000000
         when "100001100111" => A <= "000000000000000000"; -- Line 9   Column 104   Coefficient 0.00000000
         when "100001101000" => A <= "000000000000000000"; -- Line 9   Column 105   Coefficient 0.00000000
         when "100001101001" => A <= "000000000000000000"; -- Line 9   Column 106   Coefficient 0.00000000
         when "100001101010" => A <= "000000000000000000"; -- Line 9   Column 107   Coefficient 0.00000000
         when "100001101011" => A <= "000000000000000000"; -- Line 9   Column 108   Coefficient 0.00000000
         when "100001101100" => A <= "000000000000000000"; -- Line 9   Column 109   Coefficient 0.00000000
         when "100001101101" => A <= "000000000000000000"; -- Line 9   Column 110   Coefficient 0.00000000
         when "100001101110" => A <= "000000000000000000"; -- Line 9   Column 111   Coefficient 0.00000000
         when "100001101111" => A <= "000000000000000000"; -- Line 9   Column 112   Coefficient 0.00000000
         when "100001110000" => A <= "000000000000000000"; -- Line 9   Column 113   Coefficient 0.00000000
         when "100001110001" => A <= "000000000000000000"; -- Line 9   Column 114   Coefficient 0.00000000
         when "100001110010" => A <= "000000000000000000"; -- Line 9   Column 115   Coefficient 0.00000000
         when "100001110011" => A <= "000000000000000000"; -- Line 9   Column 116   Coefficient 0.00000000
         when "100001110100" => A <= "000000000000000000"; -- Line 9   Column 117   Coefficient 0.00000000
         when "100001110101" => A <= "000000000000000000"; -- Line 9   Column 118   Coefficient 0.00000000
         when "100001110110" => A <= "000000000000000000"; -- Line 9   Column 119   Coefficient 0.00000000
         when "100001110111" => A <= "000000000000000000"; -- Line 9   Column 120   Coefficient 0.00000000
         when "100001111000" => A <= "000000000000000000"; -- Line 9   Column 121   Coefficient 0.00000000
         when "100001111001" => A <= "000000000000000000"; -- Line 9   Column 122   Coefficient 0.00000000
         when "100001111010" => A <= "000000000000000000"; -- Line 9   Column 123   Coefficient 0.00000000
         when "100001111011" => A <= "000000000000000000"; -- Line 9   Column 124   Coefficient 0.00000000
         when "100001111100" => A <= "000000000000000000"; -- Line 9   Column 125   Coefficient 0.00000000
         when "100001111101" => A <= "000000000000000000"; -- Line 9   Column 126   Coefficient 0.00000000
         when "100001111110" => A <= "000000000000000000"; -- Line 9   Column 127   Coefficient 0.00000000
         when "100001111111" => A <= "000000000000000000"; -- Line 9   Column 128   Coefficient 0.00000000
         when "100010000000" => A <= "000000000000001001"; -- Line 9   Column 129   Coefficient 0.00003433
         when "100010000001" => A <= "000000000000000011"; -- Line 9   Column 130   Coefficient 0.00001144
         when "100010000010" => A <= "111111111111001011"; -- Line 9   Column 131   Coefficient -0.00020218
         when "100010000011" => A <= "111111111110100110"; -- Line 9   Column 132   Coefficient -0.00034332
         when "100010000100" => A <= "111111111110010010"; -- Line 9   Column 133   Coefficient -0.00041962
         when "100010000101" => A <= "111111111111010011"; -- Line 9   Column 134   Coefficient -0.00017166
         when "100010000110" => A <= "000000000011111000"; -- Line 9   Column 135   Coefficient 0.00094604
         when "100010000111" => A <= "000000001000010011"; -- Line 9   Column 136   Coefficient 0.00202560
         when "100010001000" => A <= "000000001010110110"; -- Line 9   Column 137   Coefficient 0.00264740
         when "100010001001" => A <= "000000001101001100"; -- Line 9   Column 138   Coefficient 0.00321960
         when "100010001010" => A <= "000000001111111100"; -- Line 9   Column 139   Coefficient 0.00389099
         when "100010001011" => A <= "000000010000011000"; -- Line 9   Column 140   Coefficient 0.00399780
         when "100010001100" => A <= "000000001111000010"; -- Line 9   Column 141   Coefficient 0.00366974
         when "100010001101" => A <= "000000000111011010"; -- Line 9   Column 142   Coefficient 0.00180817
         when "100010001110" => A <= "111111110001010101"; -- Line 9   Column 143   Coefficient -0.00358200
         when "100010001111" => A <= "111111011001111001"; -- Line 9   Column 144   Coefficient -0.00930405
         when "100010010000" => A <= "111111000100111001"; -- Line 9   Column 145   Coefficient -0.01443100
         when "100010010001" => A <= "111110110001100001"; -- Line 9   Column 146   Coefficient -0.01916122
         when "100010010010" => A <= "111110100110010011"; -- Line 9   Column 147   Coefficient -0.02190018
         when "100010010011" => A <= "111110011011111010"; -- Line 9   Column 148   Coefficient -0.02443695
         when "100010010100" => A <= "111110010000110000"; -- Line 9   Column 149   Coefficient -0.02716064
         when "100010010101" => A <= "111110000101010011"; -- Line 9   Column 150   Coefficient -0.02995682
         when "100010010110" => A <= "111101110100001010"; -- Line 9   Column 151   Coefficient -0.03414154
         when "100010010111" => A <= "111101100110110000"; -- Line 9   Column 152   Coefficient -0.03741455
         when "100010011000" => A <= "111101100010101111"; -- Line 9   Column 153   Coefficient -0.03839493
         when "100010011001" => A <= "111101100010001110"; -- Line 9   Column 154   Coefficient -0.03852081
         when "100010011010" => A <= "111101100000101101"; -- Line 9   Column 155   Coefficient -0.03889084
         when "100010011011" => A <= "111101101011101110"; -- Line 9   Column 156   Coefficient -0.03620148
         when "100010011100" => A <= "111110000010011110"; -- Line 9   Column 157   Coefficient -0.03064728
         when "100010011101" => A <= "111110110101100100"; -- Line 9   Column 158   Coefficient -0.01817322
         when "100010011110" => A <= "000000100101011001"; -- Line 9   Column 159   Coefficient 0.00912857
         when "100010011111" => A <= "000010011110111100"; -- Line 9   Column 160   Coefficient 0.03880310
         when "100010100000" => A <= "000100010010000101"; -- Line 9   Column 161   Coefficient 0.06691360
         when "100010100001" => A <= "000110000101110011"; -- Line 9   Column 162   Coefficient 0.09516525
         when "100010100010" => A <= "000111100110110001"; -- Line 9   Column 163   Coefficient 0.11883926
         when "100010100011" => A <= "001001000110101001"; -- Line 9   Column 164   Coefficient 0.14224625
         when "100010100100" => A <= "001010101100000111"; -- Line 9   Column 165   Coefficient 0.16701889
         when "100010100101" => A <= "001100001011101000"; -- Line 9   Column 166   Coefficient 0.19033813
         when "100010100110" => A <= "001101100011111111"; -- Line 9   Column 167   Coefficient 0.21191025
         when "100010100111" => A <= "001110110101010100"; -- Line 9   Column 168   Coefficient 0.23176575
         when "100010101000" => A <= "001111111010100001"; -- Line 9   Column 169   Coefficient 0.24866104
         when "100010101001" => A <= "010000111010100101"; -- Line 9   Column 170   Coefficient 0.26430130
         when "100010101010" => A <= "010010000001100011"; -- Line 9   Column 171   Coefficient 0.28162766
         when "100010101011" => A <= "010010110100110100"; -- Line 9   Column 172   Coefficient 0.29414368
         when "100010101100" => A <= "010011010010100110"; -- Line 9   Column 173   Coefficient 0.30141449
         when "100010101101" => A <= "010011000101100111"; -- Line 9   Column 174   Coefficient 0.29824448
         when "100010101110" => A <= "010001011110001011"; -- Line 9   Column 175   Coefficient 0.27299118
         when "100010101111" => A <= "001111100101110011"; -- Line 9   Column 176   Coefficient 0.24360275
         when "100010110000" => A <= "001101110100101001"; -- Line 9   Column 177   Coefficient 0.21597672
         when "100010110001" => A <= "001011111101111010"; -- Line 9   Column 178   Coefficient 0.18698883
         when "100010110010" => A <= "001010011001111000"; -- Line 9   Column 179   Coefficient 0.16256714
         when "100010110011" => A <= "001000110101000000"; -- Line 9   Column 180   Coefficient 0.13793945
         when "100010110100" => A <= "000111000101010101"; -- Line 9   Column 181   Coefficient 0.11067581
         when "100010110101" => A <= "000101100000010101"; -- Line 9   Column 182   Coefficient 0.08601761
         when "100010110110" => A <= "000100010011001101"; -- Line 9   Column 183   Coefficient 0.06718826
         when "100010110111" => A <= "000011001010010011"; -- Line 9   Column 184   Coefficient 0.04938889
         when "100010111000" => A <= "000010000100001011"; -- Line 9   Column 185   Coefficient 0.03226852
         when "100010111001" => A <= "000000111110100110"; -- Line 9   Column 186   Coefficient 0.01528168
         when "100010111010" => A <= "111111101010001000"; -- Line 9   Column 187   Coefficient -0.00534058
         when "100010111011" => A <= "111110100000101100"; -- Line 9   Column 188   Coefficient -0.02326965
         when "100010111100" => A <= "111101100111001110"; -- Line 9   Column 189   Coefficient -0.03730011
         when "100010111101" => A <= "111101000110110001"; -- Line 9   Column 190   Coefficient -0.04522324
         when "100010111110" => A <= "111101011101101101"; -- Line 9   Column 191   Coefficient -0.03962326
         when "100010111111" => A <= "111101111110110001"; -- Line 9   Column 192   Coefficient -0.03155136
         when "100011000000" => A <= "111110011010010101"; -- Line 9   Column 193   Coefficient -0.02482224
         when "100011000001" => A <= "111110111010000001"; -- Line 9   Column 194   Coefficient -0.01708603
         when "100011000010" => A <= "111111010000101110"; -- Line 9   Column 195   Coefficient -0.01154327
         when "100011000011" => A <= "111111100111100010"; -- Line 9   Column 196   Coefficient -0.00597382
         when "100011000100" => A <= "000000000100100100"; -- Line 9   Column 197   Coefficient 0.00111389
         when "100011000101" => A <= "000000011000110111"; -- Line 9   Column 198   Coefficient 0.00606918
         when "100011000110" => A <= "000000010111101010"; -- Line 9   Column 199   Coefficient 0.00577545
         when "100011000111" => A <= "000000010100111001"; -- Line 9   Column 200   Coefficient 0.00510025
         when "100011001000" => A <= "000000010100110111"; -- Line 9   Column 201   Coefficient 0.00509262
         when "100011001001" => A <= "000000010110010000"; -- Line 9   Column 202   Coefficient 0.00543213
         when "100011001010" => A <= "000000100010100100"; -- Line 9   Column 203   Coefficient 0.00843811
         when "100011001011" => A <= "000000101101010111"; -- Line 9   Column 204   Coefficient 0.01107407
         when "100011001100" => A <= "000000110010101110"; -- Line 9   Column 205   Coefficient 0.01238251
         when "100011001101" => A <= "000000110100010110"; -- Line 9   Column 206   Coefficient 0.01277924
         when "100011001110" => A <= "000000101011110101"; -- Line 9   Column 207   Coefficient 0.01070023
         when "100011001111" => A <= "000000100001110011"; -- Line 9   Column 208   Coefficient 0.00825119
         when "100011010000" => A <= "000000011001110100"; -- Line 9   Column 209   Coefficient 0.00630188
         when "100011010001" => A <= "000000010001001000"; -- Line 9   Column 210   Coefficient 0.00418091
         when "100011010010" => A <= "000000001001011000"; -- Line 9   Column 211   Coefficient 0.00228882
         when "100011010011" => A <= "000000000010010011"; -- Line 9   Column 212   Coefficient 0.00056076
         when "100011010100" => A <= "111111111010111001"; -- Line 9   Column 213   Coefficient -0.00124741
         when "100011010101" => A <= "111111110110011111"; -- Line 9   Column 214   Coefficient -0.00232315
         when "100011010110" => A <= "111111111001000110"; -- Line 9   Column 215   Coefficient -0.00168610
         when "100011010111" => A <= "111111111100011110"; -- Line 9   Column 216   Coefficient -0.00086212
         when "100011011000" => A <= "111111111110110111"; -- Line 9   Column 217   Coefficient -0.00027847
         when "100011011001" => A <= "000000000001001011"; -- Line 9   Column 218   Coefficient 0.00028610
         when "100011011010" => A <= "000000000001001000"; -- Line 9   Column 219   Coefficient 0.00027466
         when "100011011011" => A <= "000000000001000010"; -- Line 9   Column 220   Coefficient 0.00025177
         when "100011011100" => A <= "000000000001111110"; -- Line 9   Column 221   Coefficient 0.00048065
         when "100011011101" => A <= "000000000010010101"; -- Line 9   Column 222   Coefficient 0.00056839
         when "100011011110" => A <= "000000000001100101"; -- Line 9   Column 223   Coefficient 0.00038528
         when "100011011111" => A <= "000000000000110011"; -- Line 9   Column 224   Coefficient 0.00019455
         when "100011100000" => A <= "000000000000000111"; -- Line 9   Column 225   Coefficient 0.00002670
         when "100011100001" => A <= "111111111111100110"; -- Line 9   Column 226   Coefficient -0.00009918
         when "100011100010" => A <= "111111111111110100"; -- Line 9   Column 227   Coefficient -0.00004578
         when "100011100011" => A <= "000000000000000011"; -- Line 9   Column 228   Coefficient 0.00001144
         when "100011100100" => A <= "000000000000000100"; -- Line 9   Column 229   Coefficient 0.00001526
         when "100011100101" => A <= "000000000000000110"; -- Line 9   Column 230   Coefficient 0.00002289
         when "100011100110" => A <= "000000000000000011"; -- Line 9   Column 231   Coefficient 0.00001144
         when "100011100111" => A <= "111111111111111111"; -- Line 9   Column 232   Coefficient -0.00000381
         when "100011101000" => A <= "000000000000000000"; -- Line 9   Column 233   Coefficient 0.00000000
         when "100011101001" => A <= "000000000000000000"; -- Line 9   Column 234   Coefficient 0.00000000
         when "100011101010" => A <= "000000000000000000"; -- Line 9   Column 235   Coefficient 0.00000000
         when "100011101011" => A <= "000000000000000000"; -- Line 9   Column 236   Coefficient 0.00000000
         when "100011101100" => A <= "000000000000000000"; -- Line 9   Column 237   Coefficient 0.00000000
         when "100011101101" => A <= "000000000000000000"; -- Line 9   Column 238   Coefficient 0.00000000
         when "100011101110" => A <= "000000000000000000"; -- Line 9   Column 239   Coefficient 0.00000000
         when "100011101111" => A <= "000000000000000000"; -- Line 9   Column 240   Coefficient 0.00000000
         when "100011110000" => A <= "000000000000000000"; -- Line 9   Column 241   Coefficient 0.00000000
         when "100011110001" => A <= "000000000000000000"; -- Line 9   Column 242   Coefficient 0.00000000
         when "100011110010" => A <= "000000000000000000"; -- Line 9   Column 243   Coefficient 0.00000000
         when "100011110011" => A <= "000000000000000000"; -- Line 9   Column 244   Coefficient 0.00000000
         when "100011110100" => A <= "000000000000000000"; -- Line 9   Column 245   Coefficient 0.00000000
         when "100011110101" => A <= "000000000000000000"; -- Line 9   Column 246   Coefficient 0.00000000
         when "100011110110" => A <= "000000000000000000"; -- Line 9   Column 247   Coefficient 0.00000000
         when "100011110111" => A <= "000000000000000000"; -- Line 9   Column 248   Coefficient 0.00000000
         when "100011111000" => A <= "000000000000000000"; -- Line 9   Column 249   Coefficient 0.00000000
         when "100011111001" => A <= "000000000000000000"; -- Line 9   Column 250   Coefficient 0.00000000
         when "100011111010" => A <= "000000000000000000"; -- Line 9   Column 251   Coefficient 0.00000000
         when "100011111011" => A <= "000000000000000000"; -- Line 9   Column 252   Coefficient 0.00000000
         when "100011111100" => A <= "000000000000000000"; -- Line 9   Column 253   Coefficient 0.00000000
         when "100011111101" => A <= "000000000000000000"; -- Line 9   Column 254   Coefficient 0.00000000
         when "100011111110" => A <= "000000000000000000"; -- Line 9   Column 255   Coefficient 0.00000000
         when "100011111111" => A <= "000000000000000000"; -- Line 9   Column 256   Coefficient 0.00000000
         when "100100000000" => A <= "000000000000000000"; -- Line 10   Column 1   Coefficient 0.00000000
         when "100100000001" => A <= "000000000000000000"; -- Line 10   Column 2   Coefficient 0.00000000
         when "100100000010" => A <= "000000000000000000"; -- Line 10   Column 3   Coefficient 0.00000000
         when "100100000011" => A <= "000000000000000000"; -- Line 10   Column 4   Coefficient 0.00000000
         when "100100000100" => A <= "000000000000000000"; -- Line 10   Column 5   Coefficient 0.00000000
         when "100100000101" => A <= "000000000000000000"; -- Line 10   Column 6   Coefficient 0.00000000
         when "100100000110" => A <= "000000000000000000"; -- Line 10   Column 7   Coefficient 0.00000000
         when "100100000111" => A <= "000000000000000000"; -- Line 10   Column 8   Coefficient 0.00000000
         when "100100001000" => A <= "000000000000000000"; -- Line 10   Column 9   Coefficient 0.00000000
         when "100100001001" => A <= "000000000000000000"; -- Line 10   Column 10   Coefficient 0.00000000
         when "100100001010" => A <= "000000000000000000"; -- Line 10   Column 11   Coefficient 0.00000000
         when "100100001011" => A <= "000000000000000000"; -- Line 10   Column 12   Coefficient 0.00000000
         when "100100001100" => A <= "000000000000000000"; -- Line 10   Column 13   Coefficient 0.00000000
         when "100100001101" => A <= "000000000000000000"; -- Line 10   Column 14   Coefficient 0.00000000
         when "100100001110" => A <= "000000000000000000"; -- Line 10   Column 15   Coefficient 0.00000000
         when "100100001111" => A <= "000000000000000000"; -- Line 10   Column 16   Coefficient 0.00000000
         when "100100010000" => A <= "000000000000000000"; -- Line 10   Column 17   Coefficient 0.00000000
         when "100100010001" => A <= "000000000000000000"; -- Line 10   Column 18   Coefficient 0.00000000
         when "100100010010" => A <= "000000000000000000"; -- Line 10   Column 19   Coefficient 0.00000000
         when "100100010011" => A <= "000000000000000000"; -- Line 10   Column 20   Coefficient 0.00000000
         when "100100010100" => A <= "000000000000000000"; -- Line 10   Column 21   Coefficient 0.00000000
         when "100100010101" => A <= "000000000000000000"; -- Line 10   Column 22   Coefficient 0.00000000
         when "100100010110" => A <= "000000000000000000"; -- Line 10   Column 23   Coefficient 0.00000000
         when "100100010111" => A <= "000000000000000000"; -- Line 10   Column 24   Coefficient 0.00000000
         when "100100011000" => A <= "000000000000000000"; -- Line 10   Column 25   Coefficient 0.00000000
         when "100100011001" => A <= "000000000000000000"; -- Line 10   Column 26   Coefficient 0.00000000
         when "100100011010" => A <= "000000000000000000"; -- Line 10   Column 27   Coefficient 0.00000000
         when "100100011011" => A <= "000000000000000000"; -- Line 10   Column 28   Coefficient 0.00000000
         when "100100011100" => A <= "000000000000000000"; -- Line 10   Column 29   Coefficient 0.00000000
         when "100100011101" => A <= "000000000000000000"; -- Line 10   Column 30   Coefficient 0.00000000
         when "100100011110" => A <= "000000000000000000"; -- Line 10   Column 31   Coefficient 0.00000000
         when "100100011111" => A <= "000000000000000000"; -- Line 10   Column 32   Coefficient 0.00000000
         when "100100100000" => A <= "000000000000000000"; -- Line 10   Column 33   Coefficient 0.00000000
         when "100100100001" => A <= "000000000000000000"; -- Line 10   Column 34   Coefficient 0.00000000
         when "100100100010" => A <= "000000000000000000"; -- Line 10   Column 35   Coefficient 0.00000000
         when "100100100011" => A <= "000000000000000000"; -- Line 10   Column 36   Coefficient 0.00000000
         when "100100100100" => A <= "000000000000000000"; -- Line 10   Column 37   Coefficient 0.00000000
         when "100100100101" => A <= "000000000000000000"; -- Line 10   Column 38   Coefficient 0.00000000
         when "100100100110" => A <= "000000000000000000"; -- Line 10   Column 39   Coefficient 0.00000000
         when "100100100111" => A <= "000000000000000000"; -- Line 10   Column 40   Coefficient 0.00000000
         when "100100101000" => A <= "000000000000000000"; -- Line 10   Column 41   Coefficient 0.00000000
         when "100100101001" => A <= "000000000000000000"; -- Line 10   Column 42   Coefficient 0.00000000
         when "100100101010" => A <= "000000000000000000"; -- Line 10   Column 43   Coefficient 0.00000000
         when "100100101011" => A <= "000000000000000000"; -- Line 10   Column 44   Coefficient 0.00000000
         when "100100101100" => A <= "000000000000000000"; -- Line 10   Column 45   Coefficient 0.00000000
         when "100100101101" => A <= "000000000000000000"; -- Line 10   Column 46   Coefficient 0.00000000
         when "100100101110" => A <= "000000000000000000"; -- Line 10   Column 47   Coefficient 0.00000000
         when "100100101111" => A <= "000000000000000000"; -- Line 10   Column 48   Coefficient 0.00000000
         when "100100110000" => A <= "000000000000000000"; -- Line 10   Column 49   Coefficient 0.00000000
         when "100100110001" => A <= "000000000000000000"; -- Line 10   Column 50   Coefficient 0.00000000
         when "100100110010" => A <= "000000000000000000"; -- Line 10   Column 51   Coefficient 0.00000000
         when "100100110011" => A <= "000000000000000000"; -- Line 10   Column 52   Coefficient 0.00000000
         when "100100110100" => A <= "000000000000000000"; -- Line 10   Column 53   Coefficient 0.00000000
         when "100100110101" => A <= "000000000000000000"; -- Line 10   Column 54   Coefficient 0.00000000
         when "100100110110" => A <= "000000000000000000"; -- Line 10   Column 55   Coefficient 0.00000000
         when "100100110111" => A <= "000000000000000000"; -- Line 10   Column 56   Coefficient 0.00000000
         when "100100111000" => A <= "000000000000000000"; -- Line 10   Column 57   Coefficient 0.00000000
         when "100100111001" => A <= "000000000000000000"; -- Line 10   Column 58   Coefficient 0.00000000
         when "100100111010" => A <= "000000000000000000"; -- Line 10   Column 59   Coefficient 0.00000000
         when "100100111011" => A <= "000000000000000000"; -- Line 10   Column 60   Coefficient 0.00000000
         when "100100111100" => A <= "000000000000000000"; -- Line 10   Column 61   Coefficient 0.00000000
         when "100100111101" => A <= "000000000000000000"; -- Line 10   Column 62   Coefficient 0.00000000
         when "100100111110" => A <= "000000000000000000"; -- Line 10   Column 63   Coefficient 0.00000000
         when "100100111111" => A <= "000000000000000000"; -- Line 10   Column 64   Coefficient 0.00000000
         when "100101000000" => A <= "000000000000000000"; -- Line 10   Column 65   Coefficient 0.00000000
         when "100101000001" => A <= "000000000000000000"; -- Line 10   Column 66   Coefficient 0.00000000
         when "100101000010" => A <= "000000000000000000"; -- Line 10   Column 67   Coefficient 0.00000000
         when "100101000011" => A <= "000000000000000000"; -- Line 10   Column 68   Coefficient 0.00000000
         when "100101000100" => A <= "000000000000000000"; -- Line 10   Column 69   Coefficient 0.00000000
         when "100101000101" => A <= "000000000000000000"; -- Line 10   Column 70   Coefficient 0.00000000
         when "100101000110" => A <= "000000000000000000"; -- Line 10   Column 71   Coefficient 0.00000000
         when "100101000111" => A <= "000000000000000000"; -- Line 10   Column 72   Coefficient 0.00000000
         when "100101001000" => A <= "000000000000000000"; -- Line 10   Column 73   Coefficient 0.00000000
         when "100101001001" => A <= "000000000000000000"; -- Line 10   Column 74   Coefficient 0.00000000
         when "100101001010" => A <= "000000000000000000"; -- Line 10   Column 75   Coefficient 0.00000000
         when "100101001011" => A <= "000000000000000000"; -- Line 10   Column 76   Coefficient 0.00000000
         when "100101001100" => A <= "000000000000000000"; -- Line 10   Column 77   Coefficient 0.00000000
         when "100101001101" => A <= "000000000000000000"; -- Line 10   Column 78   Coefficient 0.00000000
         when "100101001110" => A <= "000000000000000000"; -- Line 10   Column 79   Coefficient 0.00000000
         when "100101001111" => A <= "000000000000000000"; -- Line 10   Column 80   Coefficient 0.00000000
         when "100101010000" => A <= "000000000000000000"; -- Line 10   Column 81   Coefficient 0.00000000
         when "100101010001" => A <= "000000000000000000"; -- Line 10   Column 82   Coefficient 0.00000000
         when "100101010010" => A <= "000000000000000000"; -- Line 10   Column 83   Coefficient 0.00000000
         when "100101010011" => A <= "000000000000000000"; -- Line 10   Column 84   Coefficient 0.00000000
         when "100101010100" => A <= "000000000000000000"; -- Line 10   Column 85   Coefficient 0.00000000
         when "100101010101" => A <= "000000000000000000"; -- Line 10   Column 86   Coefficient 0.00000000
         when "100101010110" => A <= "000000000000000000"; -- Line 10   Column 87   Coefficient 0.00000000
         when "100101010111" => A <= "000000000000000000"; -- Line 10   Column 88   Coefficient 0.00000000
         when "100101011000" => A <= "000000000000000000"; -- Line 10   Column 89   Coefficient 0.00000000
         when "100101011001" => A <= "000000000000000000"; -- Line 10   Column 90   Coefficient 0.00000000
         when "100101011010" => A <= "000000000000000000"; -- Line 10   Column 91   Coefficient 0.00000000
         when "100101011011" => A <= "000000000000000000"; -- Line 10   Column 92   Coefficient 0.00000000
         when "100101011100" => A <= "000000000000000000"; -- Line 10   Column 93   Coefficient 0.00000000
         when "100101011101" => A <= "000000000000000000"; -- Line 10   Column 94   Coefficient 0.00000000
         when "100101011110" => A <= "000000000000000000"; -- Line 10   Column 95   Coefficient 0.00000000
         when "100101011111" => A <= "000000000000000000"; -- Line 10   Column 96   Coefficient 0.00000000
         when "100101100000" => A <= "000000000000000000"; -- Line 10   Column 97   Coefficient 0.00000000
         when "100101100001" => A <= "000000000000000000"; -- Line 10   Column 98   Coefficient 0.00000000
         when "100101100010" => A <= "000000000000000000"; -- Line 10   Column 99   Coefficient 0.00000000
         when "100101100011" => A <= "000000000000000000"; -- Line 10   Column 100   Coefficient 0.00000000
         when "100101100100" => A <= "000000000000000000"; -- Line 10   Column 101   Coefficient 0.00000000
         when "100101100101" => A <= "000000000000000000"; -- Line 10   Column 102   Coefficient 0.00000000
         when "100101100110" => A <= "000000000000000000"; -- Line 10   Column 103   Coefficient 0.00000000
         when "100101100111" => A <= "000000000000000000"; -- Line 10   Column 104   Coefficient 0.00000000
         when "100101101000" => A <= "000000000000000000"; -- Line 10   Column 105   Coefficient 0.00000000
         when "100101101001" => A <= "000000000000000000"; -- Line 10   Column 106   Coefficient 0.00000000
         when "100101101010" => A <= "000000000000000000"; -- Line 10   Column 107   Coefficient 0.00000000
         when "100101101011" => A <= "000000000000000000"; -- Line 10   Column 108   Coefficient 0.00000000
         when "100101101100" => A <= "000000000000000000"; -- Line 10   Column 109   Coefficient 0.00000000
         when "100101101101" => A <= "000000000000000000"; -- Line 10   Column 110   Coefficient 0.00000000
         when "100101101110" => A <= "000000000000000000"; -- Line 10   Column 111   Coefficient 0.00000000
         when "100101101111" => A <= "000000000000000000"; -- Line 10   Column 112   Coefficient 0.00000000
         when "100101110000" => A <= "000000000000000000"; -- Line 10   Column 113   Coefficient 0.00000000
         when "100101110001" => A <= "000000000000000000"; -- Line 10   Column 114   Coefficient 0.00000000
         when "100101110010" => A <= "000000000000000000"; -- Line 10   Column 115   Coefficient 0.00000000
         when "100101110011" => A <= "000000000000000000"; -- Line 10   Column 116   Coefficient 0.00000000
         when "100101110100" => A <= "000000000000000000"; -- Line 10   Column 117   Coefficient 0.00000000
         when "100101110101" => A <= "000000000000000000"; -- Line 10   Column 118   Coefficient 0.00000000
         when "100101110110" => A <= "000000000000000000"; -- Line 10   Column 119   Coefficient 0.00000000
         when "100101110111" => A <= "000000000000000000"; -- Line 10   Column 120   Coefficient 0.00000000
         when "100101111000" => A <= "000000000000000000"; -- Line 10   Column 121   Coefficient 0.00000000
         when "100101111001" => A <= "000000000000000000"; -- Line 10   Column 122   Coefficient 0.00000000
         when "100101111010" => A <= "000000000000000000"; -- Line 10   Column 123   Coefficient 0.00000000
         when "100101111011" => A <= "000000000000000000"; -- Line 10   Column 124   Coefficient 0.00000000
         when "100101111100" => A <= "000000000000000000"; -- Line 10   Column 125   Coefficient 0.00000000
         when "100101111101" => A <= "000000000000000000"; -- Line 10   Column 126   Coefficient 0.00000000
         when "100101111110" => A <= "000000000000000000"; -- Line 10   Column 127   Coefficient 0.00000000
         when "100101111111" => A <= "000000000000000000"; -- Line 10   Column 128   Coefficient 0.00000000
         when "100110000000" => A <= "000000000000000000"; -- Line 10   Column 129   Coefficient 0.00000000
         when "100110000001" => A <= "000000000000000000"; -- Line 10   Column 130   Coefficient 0.00000000
         when "100110000010" => A <= "000000000000000000"; -- Line 10   Column 131   Coefficient 0.00000000
         when "100110000011" => A <= "000000000000000000"; -- Line 10   Column 132   Coefficient 0.00000000
         when "100110000100" => A <= "000000000000000000"; -- Line 10   Column 133   Coefficient 0.00000000
         when "100110000101" => A <= "000000000000000000"; -- Line 10   Column 134   Coefficient 0.00000000
         when "100110000110" => A <= "000000000000000000"; -- Line 10   Column 135   Coefficient 0.00000000
         when "100110000111" => A <= "000000000000000000"; -- Line 10   Column 136   Coefficient 0.00000000
         when "100110001000" => A <= "000000000000000000"; -- Line 10   Column 137   Coefficient 0.00000000
         when "100110001001" => A <= "000000000000000000"; -- Line 10   Column 138   Coefficient 0.00000000
         when "100110001010" => A <= "000000000000000000"; -- Line 10   Column 139   Coefficient 0.00000000
         when "100110001011" => A <= "000000000000000000"; -- Line 10   Column 140   Coefficient 0.00000000
         when "100110001100" => A <= "000000000000000000"; -- Line 10   Column 141   Coefficient 0.00000000
         when "100110001101" => A <= "000000000000000000"; -- Line 10   Column 142   Coefficient 0.00000000
         when "100110001110" => A <= "000000000000000000"; -- Line 10   Column 143   Coefficient 0.00000000
         when "100110001111" => A <= "000000000000000000"; -- Line 10   Column 144   Coefficient 0.00000000
         when "100110010000" => A <= "000000000000001001"; -- Line 10   Column 145   Coefficient 0.00003433
         when "100110010001" => A <= "000000000000000011"; -- Line 10   Column 146   Coefficient 0.00001144
         when "100110010010" => A <= "111111111111001011"; -- Line 10   Column 147   Coefficient -0.00020218
         when "100110010011" => A <= "111111111110100110"; -- Line 10   Column 148   Coefficient -0.00034332
         when "100110010100" => A <= "111111111110010010"; -- Line 10   Column 149   Coefficient -0.00041962
         when "100110010101" => A <= "111111111111010011"; -- Line 10   Column 150   Coefficient -0.00017166
         when "100110010110" => A <= "000000000011111000"; -- Line 10   Column 151   Coefficient 0.00094604
         when "100110010111" => A <= "000000001000010011"; -- Line 10   Column 152   Coefficient 0.00202560
         when "100110011000" => A <= "000000001010110110"; -- Line 10   Column 153   Coefficient 0.00264740
         when "100110011001" => A <= "000000001101001100"; -- Line 10   Column 154   Coefficient 0.00321960
         when "100110011010" => A <= "000000001111111100"; -- Line 10   Column 155   Coefficient 0.00389099
         when "100110011011" => A <= "000000010000011000"; -- Line 10   Column 156   Coefficient 0.00399780
         when "100110011100" => A <= "000000001111000010"; -- Line 10   Column 157   Coefficient 0.00366974
         when "100110011101" => A <= "000000000111011010"; -- Line 10   Column 158   Coefficient 0.00180817
         when "100110011110" => A <= "111111110001010101"; -- Line 10   Column 159   Coefficient -0.00358200
         when "100110011111" => A <= "111111011001111001"; -- Line 10   Column 160   Coefficient -0.00930405
         when "100110100000" => A <= "111111000100111001"; -- Line 10   Column 161   Coefficient -0.01443100
         when "100110100001" => A <= "111110110001100001"; -- Line 10   Column 162   Coefficient -0.01916122
         when "100110100010" => A <= "111110100110010011"; -- Line 10   Column 163   Coefficient -0.02190018
         when "100110100011" => A <= "111110011011111010"; -- Line 10   Column 164   Coefficient -0.02443695
         when "100110100100" => A <= "111110010000110000"; -- Line 10   Column 165   Coefficient -0.02716064
         when "100110100101" => A <= "111110000101010011"; -- Line 10   Column 166   Coefficient -0.02995682
         when "100110100110" => A <= "111101110100001010"; -- Line 10   Column 167   Coefficient -0.03414154
         when "100110100111" => A <= "111101100110110000"; -- Line 10   Column 168   Coefficient -0.03741455
         when "100110101000" => A <= "111101100010101111"; -- Line 10   Column 169   Coefficient -0.03839493
         when "100110101001" => A <= "111101100010001110"; -- Line 10   Column 170   Coefficient -0.03852081
         when "100110101010" => A <= "111101100000101101"; -- Line 10   Column 171   Coefficient -0.03889084
         when "100110101011" => A <= "111101101011101110"; -- Line 10   Column 172   Coefficient -0.03620148
         when "100110101100" => A <= "111110000010011110"; -- Line 10   Column 173   Coefficient -0.03064728
         when "100110101101" => A <= "111110110101100100"; -- Line 10   Column 174   Coefficient -0.01817322
         when "100110101110" => A <= "000000100101011001"; -- Line 10   Column 175   Coefficient 0.00912857
         when "100110101111" => A <= "000010011110111100"; -- Line 10   Column 176   Coefficient 0.03880310
         when "100110110000" => A <= "000100010010000101"; -- Line 10   Column 177   Coefficient 0.06691360
         when "100110110001" => A <= "000110000101110011"; -- Line 10   Column 178   Coefficient 0.09516525
         when "100110110010" => A <= "000111100110110001"; -- Line 10   Column 179   Coefficient 0.11883926
         when "100110110011" => A <= "001001000110101001"; -- Line 10   Column 180   Coefficient 0.14224625
         when "100110110100" => A <= "001010101100000111"; -- Line 10   Column 181   Coefficient 0.16701889
         when "100110110101" => A <= "001100001011101000"; -- Line 10   Column 182   Coefficient 0.19033813
         when "100110110110" => A <= "001101100011111111"; -- Line 10   Column 183   Coefficient 0.21191025
         when "100110110111" => A <= "001110110101010100"; -- Line 10   Column 184   Coefficient 0.23176575
         when "100110111000" => A <= "001111111010100001"; -- Line 10   Column 185   Coefficient 0.24866104
         when "100110111001" => A <= "010000111010100101"; -- Line 10   Column 186   Coefficient 0.26430130
         when "100110111010" => A <= "010010000001100011"; -- Line 10   Column 187   Coefficient 0.28162766
         when "100110111011" => A <= "010010110100110100"; -- Line 10   Column 188   Coefficient 0.29414368
         when "100110111100" => A <= "010011010010100110"; -- Line 10   Column 189   Coefficient 0.30141449
         when "100110111101" => A <= "010011000101100111"; -- Line 10   Column 190   Coefficient 0.29824448
         when "100110111110" => A <= "010001011110001011"; -- Line 10   Column 191   Coefficient 0.27299118
         when "100110111111" => A <= "001111100101110011"; -- Line 10   Column 192   Coefficient 0.24360275
         when "100111000000" => A <= "001101110100101001"; -- Line 10   Column 193   Coefficient 0.21597672
         when "100111000001" => A <= "001011111101111010"; -- Line 10   Column 194   Coefficient 0.18698883
         when "100111000010" => A <= "001010011001111000"; -- Line 10   Column 195   Coefficient 0.16256714
         when "100111000011" => A <= "001000110101000000"; -- Line 10   Column 196   Coefficient 0.13793945
         when "100111000100" => A <= "000111000101010101"; -- Line 10   Column 197   Coefficient 0.11067581
         when "100111000101" => A <= "000101100000010101"; -- Line 10   Column 198   Coefficient 0.08601761
         when "100111000110" => A <= "000100010011001101"; -- Line 10   Column 199   Coefficient 0.06718826
         when "100111000111" => A <= "000011001010010011"; -- Line 10   Column 200   Coefficient 0.04938889
         when "100111001000" => A <= "000010000100001011"; -- Line 10   Column 201   Coefficient 0.03226852
         when "100111001001" => A <= "000000111110100110"; -- Line 10   Column 202   Coefficient 0.01528168
         when "100111001010" => A <= "111111101010001000"; -- Line 10   Column 203   Coefficient -0.00534058
         when "100111001011" => A <= "111110100000101100"; -- Line 10   Column 204   Coefficient -0.02326965
         when "100111001100" => A <= "111101100111001110"; -- Line 10   Column 205   Coefficient -0.03730011
         when "100111001101" => A <= "111101000110110001"; -- Line 10   Column 206   Coefficient -0.04522324
         when "100111001110" => A <= "111101011101101101"; -- Line 10   Column 207   Coefficient -0.03962326
         when "100111001111" => A <= "111101111110110001"; -- Line 10   Column 208   Coefficient -0.03155136
         when "100111010000" => A <= "111110011010010101"; -- Line 10   Column 209   Coefficient -0.02482224
         when "100111010001" => A <= "111110111010000001"; -- Line 10   Column 210   Coefficient -0.01708603
         when "100111010010" => A <= "111111010000101110"; -- Line 10   Column 211   Coefficient -0.01154327
         when "100111010011" => A <= "111111100111100010"; -- Line 10   Column 212   Coefficient -0.00597382
         when "100111010100" => A <= "000000000100100100"; -- Line 10   Column 213   Coefficient 0.00111389
         when "100111010101" => A <= "000000011000110111"; -- Line 10   Column 214   Coefficient 0.00606918
         when "100111010110" => A <= "000000010111101010"; -- Line 10   Column 215   Coefficient 0.00577545
         when "100111010111" => A <= "000000010100111001"; -- Line 10   Column 216   Coefficient 0.00510025
         when "100111011000" => A <= "000000010100110111"; -- Line 10   Column 217   Coefficient 0.00509262
         when "100111011001" => A <= "000000010110010000"; -- Line 10   Column 218   Coefficient 0.00543213
         when "100111011010" => A <= "000000100010100100"; -- Line 10   Column 219   Coefficient 0.00843811
         when "100111011011" => A <= "000000101101010111"; -- Line 10   Column 220   Coefficient 0.01107407
         when "100111011100" => A <= "000000110010101110"; -- Line 10   Column 221   Coefficient 0.01238251
         when "100111011101" => A <= "000000110100010110"; -- Line 10   Column 222   Coefficient 0.01277924
         when "100111011110" => A <= "000000101011110101"; -- Line 10   Column 223   Coefficient 0.01070023
         when "100111011111" => A <= "000000100001110011"; -- Line 10   Column 224   Coefficient 0.00825119
         when "100111100000" => A <= "000000011001110100"; -- Line 10   Column 225   Coefficient 0.00630188
         when "100111100001" => A <= "000000010001001000"; -- Line 10   Column 226   Coefficient 0.00418091
         when "100111100010" => A <= "000000001001011000"; -- Line 10   Column 227   Coefficient 0.00228882
         when "100111100011" => A <= "000000000010010011"; -- Line 10   Column 228   Coefficient 0.00056076
         when "100111100100" => A <= "111111111010111001"; -- Line 10   Column 229   Coefficient -0.00124741
         when "100111100101" => A <= "111111110110011111"; -- Line 10   Column 230   Coefficient -0.00232315
         when "100111100110" => A <= "111111111001000110"; -- Line 10   Column 231   Coefficient -0.00168610
         when "100111100111" => A <= "111111111100011110"; -- Line 10   Column 232   Coefficient -0.00086212
         when "100111101000" => A <= "111111111110110111"; -- Line 10   Column 233   Coefficient -0.00027847
         when "100111101001" => A <= "000000000001001011"; -- Line 10   Column 234   Coefficient 0.00028610
         when "100111101010" => A <= "000000000001001000"; -- Line 10   Column 235   Coefficient 0.00027466
         when "100111101011" => A <= "000000000001000010"; -- Line 10   Column 236   Coefficient 0.00025177
         when "100111101100" => A <= "000000000001111110"; -- Line 10   Column 237   Coefficient 0.00048065
         when "100111101101" => A <= "000000000010010101"; -- Line 10   Column 238   Coefficient 0.00056839
         when "100111101110" => A <= "000000000001100101"; -- Line 10   Column 239   Coefficient 0.00038528
         when "100111101111" => A <= "000000000000110011"; -- Line 10   Column 240   Coefficient 0.00019455
         when "100111110000" => A <= "000000000000000111"; -- Line 10   Column 241   Coefficient 0.00002670
         when "100111110001" => A <= "111111111111100110"; -- Line 10   Column 242   Coefficient -0.00009918
         when "100111110010" => A <= "111111111111110100"; -- Line 10   Column 243   Coefficient -0.00004578
         when "100111110011" => A <= "000000000000000011"; -- Line 10   Column 244   Coefficient 0.00001144
         when "100111110100" => A <= "000000000000000100"; -- Line 10   Column 245   Coefficient 0.00001526
         when "100111110101" => A <= "000000000000000110"; -- Line 10   Column 246   Coefficient 0.00002289
         when "100111110110" => A <= "000000000000000011"; -- Line 10   Column 247   Coefficient 0.00001144
         when "100111110111" => A <= "111111111111111111"; -- Line 10   Column 248   Coefficient -0.00000381
         when "100111111000" => A <= "000000000000000000"; -- Line 10   Column 249   Coefficient 0.00000000
         when "100111111001" => A <= "000000000000000000"; -- Line 10   Column 250   Coefficient 0.00000000
         when "100111111010" => A <= "000000000000000000"; -- Line 10   Column 251   Coefficient 0.00000000
         when "100111111011" => A <= "000000000000000000"; -- Line 10   Column 252   Coefficient 0.00000000
         when "100111111100" => A <= "000000000000000000"; -- Line 10   Column 253   Coefficient 0.00000000
         when "100111111101" => A <= "000000000000000000"; -- Line 10   Column 254   Coefficient 0.00000000
         when "100111111110" => A <= "000000000000000000"; -- Line 10   Column 255   Coefficient 0.00000000
         when "100111111111" => A <= "000000000000000000"; -- Line 10   Column 256   Coefficient 0.00000000
         when "101000000000" => A <= "000000000000000111"; -- Line 11   Column 1   Coefficient 0.00002670
         when "101000000001" => A <= "111111111111100110"; -- Line 11   Column 2   Coefficient -0.00009918
         when "101000000010" => A <= "111111111111110100"; -- Line 11   Column 3   Coefficient -0.00004578
         when "101000000011" => A <= "000000000000000011"; -- Line 11   Column 4   Coefficient 0.00001144
         when "101000000100" => A <= "000000000000000100"; -- Line 11   Column 5   Coefficient 0.00001526
         when "101000000101" => A <= "000000000000000110"; -- Line 11   Column 6   Coefficient 0.00002289
         when "101000000110" => A <= "000000000000000011"; -- Line 11   Column 7   Coefficient 0.00001144
         when "101000000111" => A <= "111111111111111111"; -- Line 11   Column 8   Coefficient -0.00000381
         when "101000001000" => A <= "000000000000000000"; -- Line 11   Column 9   Coefficient 0.00000000
         when "101000001001" => A <= "000000000000000000"; -- Line 11   Column 10   Coefficient 0.00000000
         when "101000001010" => A <= "000000000000000000"; -- Line 11   Column 11   Coefficient 0.00000000
         when "101000001011" => A <= "000000000000000000"; -- Line 11   Column 12   Coefficient 0.00000000
         when "101000001100" => A <= "000000000000000000"; -- Line 11   Column 13   Coefficient 0.00000000
         when "101000001101" => A <= "000000000000000000"; -- Line 11   Column 14   Coefficient 0.00000000
         when "101000001110" => A <= "000000000000000000"; -- Line 11   Column 15   Coefficient 0.00000000
         when "101000001111" => A <= "000000000000000000"; -- Line 11   Column 16   Coefficient 0.00000000
         when "101000010000" => A <= "000000000000000000"; -- Line 11   Column 17   Coefficient 0.00000000
         when "101000010001" => A <= "000000000000000000"; -- Line 11   Column 18   Coefficient 0.00000000
         when "101000010010" => A <= "000000000000000000"; -- Line 11   Column 19   Coefficient 0.00000000
         when "101000010011" => A <= "000000000000000000"; -- Line 11   Column 20   Coefficient 0.00000000
         when "101000010100" => A <= "000000000000000000"; -- Line 11   Column 21   Coefficient 0.00000000
         when "101000010101" => A <= "000000000000000000"; -- Line 11   Column 22   Coefficient 0.00000000
         when "101000010110" => A <= "000000000000000000"; -- Line 11   Column 23   Coefficient 0.00000000
         when "101000010111" => A <= "000000000000000000"; -- Line 11   Column 24   Coefficient 0.00000000
         when "101000011000" => A <= "000000000000000000"; -- Line 11   Column 25   Coefficient 0.00000000
         when "101000011001" => A <= "000000000000000000"; -- Line 11   Column 26   Coefficient 0.00000000
         when "101000011010" => A <= "000000000000000000"; -- Line 11   Column 27   Coefficient 0.00000000
         when "101000011011" => A <= "000000000000000000"; -- Line 11   Column 28   Coefficient 0.00000000
         when "101000011100" => A <= "000000000000000000"; -- Line 11   Column 29   Coefficient 0.00000000
         when "101000011101" => A <= "000000000000000000"; -- Line 11   Column 30   Coefficient 0.00000000
         when "101000011110" => A <= "000000000000000000"; -- Line 11   Column 31   Coefficient 0.00000000
         when "101000011111" => A <= "000000000000000000"; -- Line 11   Column 32   Coefficient 0.00000000
         when "101000100000" => A <= "000000000000000000"; -- Line 11   Column 33   Coefficient 0.00000000
         when "101000100001" => A <= "000000000000000000"; -- Line 11   Column 34   Coefficient 0.00000000
         when "101000100010" => A <= "000000000000000000"; -- Line 11   Column 35   Coefficient 0.00000000
         when "101000100011" => A <= "000000000000000000"; -- Line 11   Column 36   Coefficient 0.00000000
         when "101000100100" => A <= "000000000000000000"; -- Line 11   Column 37   Coefficient 0.00000000
         when "101000100101" => A <= "000000000000000000"; -- Line 11   Column 38   Coefficient 0.00000000
         when "101000100110" => A <= "000000000000000000"; -- Line 11   Column 39   Coefficient 0.00000000
         when "101000100111" => A <= "000000000000000000"; -- Line 11   Column 40   Coefficient 0.00000000
         when "101000101000" => A <= "000000000000000000"; -- Line 11   Column 41   Coefficient 0.00000000
         when "101000101001" => A <= "000000000000000000"; -- Line 11   Column 42   Coefficient 0.00000000
         when "101000101010" => A <= "000000000000000000"; -- Line 11   Column 43   Coefficient 0.00000000
         when "101000101011" => A <= "000000000000000000"; -- Line 11   Column 44   Coefficient 0.00000000
         when "101000101100" => A <= "000000000000000000"; -- Line 11   Column 45   Coefficient 0.00000000
         when "101000101101" => A <= "000000000000000000"; -- Line 11   Column 46   Coefficient 0.00000000
         when "101000101110" => A <= "000000000000000000"; -- Line 11   Column 47   Coefficient 0.00000000
         when "101000101111" => A <= "000000000000000000"; -- Line 11   Column 48   Coefficient 0.00000000
         when "101000110000" => A <= "000000000000000000"; -- Line 11   Column 49   Coefficient 0.00000000
         when "101000110001" => A <= "000000000000000000"; -- Line 11   Column 50   Coefficient 0.00000000
         when "101000110010" => A <= "000000000000000000"; -- Line 11   Column 51   Coefficient 0.00000000
         when "101000110011" => A <= "000000000000000000"; -- Line 11   Column 52   Coefficient 0.00000000
         when "101000110100" => A <= "000000000000000000"; -- Line 11   Column 53   Coefficient 0.00000000
         when "101000110101" => A <= "000000000000000000"; -- Line 11   Column 54   Coefficient 0.00000000
         when "101000110110" => A <= "000000000000000000"; -- Line 11   Column 55   Coefficient 0.00000000
         when "101000110111" => A <= "000000000000000000"; -- Line 11   Column 56   Coefficient 0.00000000
         when "101000111000" => A <= "000000000000000000"; -- Line 11   Column 57   Coefficient 0.00000000
         when "101000111001" => A <= "000000000000000000"; -- Line 11   Column 58   Coefficient 0.00000000
         when "101000111010" => A <= "000000000000000000"; -- Line 11   Column 59   Coefficient 0.00000000
         when "101000111011" => A <= "000000000000000000"; -- Line 11   Column 60   Coefficient 0.00000000
         when "101000111100" => A <= "000000000000000000"; -- Line 11   Column 61   Coefficient 0.00000000
         when "101000111101" => A <= "000000000000000000"; -- Line 11   Column 62   Coefficient 0.00000000
         when "101000111110" => A <= "000000000000000000"; -- Line 11   Column 63   Coefficient 0.00000000
         when "101000111111" => A <= "000000000000000000"; -- Line 11   Column 64   Coefficient 0.00000000
         when "101001000000" => A <= "000000000000000000"; -- Line 11   Column 65   Coefficient 0.00000000
         when "101001000001" => A <= "000000000000000000"; -- Line 11   Column 66   Coefficient 0.00000000
         when "101001000010" => A <= "000000000000000000"; -- Line 11   Column 67   Coefficient 0.00000000
         when "101001000011" => A <= "000000000000000000"; -- Line 11   Column 68   Coefficient 0.00000000
         when "101001000100" => A <= "000000000000000000"; -- Line 11   Column 69   Coefficient 0.00000000
         when "101001000101" => A <= "000000000000000000"; -- Line 11   Column 70   Coefficient 0.00000000
         when "101001000110" => A <= "000000000000000000"; -- Line 11   Column 71   Coefficient 0.00000000
         when "101001000111" => A <= "000000000000000000"; -- Line 11   Column 72   Coefficient 0.00000000
         when "101001001000" => A <= "000000000000000000"; -- Line 11   Column 73   Coefficient 0.00000000
         when "101001001001" => A <= "000000000000000000"; -- Line 11   Column 74   Coefficient 0.00000000
         when "101001001010" => A <= "000000000000000000"; -- Line 11   Column 75   Coefficient 0.00000000
         when "101001001011" => A <= "000000000000000000"; -- Line 11   Column 76   Coefficient 0.00000000
         when "101001001100" => A <= "000000000000000000"; -- Line 11   Column 77   Coefficient 0.00000000
         when "101001001101" => A <= "000000000000000000"; -- Line 11   Column 78   Coefficient 0.00000000
         when "101001001110" => A <= "000000000000000000"; -- Line 11   Column 79   Coefficient 0.00000000
         when "101001001111" => A <= "000000000000000000"; -- Line 11   Column 80   Coefficient 0.00000000
         when "101001010000" => A <= "000000000000000000"; -- Line 11   Column 81   Coefficient 0.00000000
         when "101001010001" => A <= "000000000000000000"; -- Line 11   Column 82   Coefficient 0.00000000
         when "101001010010" => A <= "000000000000000000"; -- Line 11   Column 83   Coefficient 0.00000000
         when "101001010011" => A <= "000000000000000000"; -- Line 11   Column 84   Coefficient 0.00000000
         when "101001010100" => A <= "000000000000000000"; -- Line 11   Column 85   Coefficient 0.00000000
         when "101001010101" => A <= "000000000000000000"; -- Line 11   Column 86   Coefficient 0.00000000
         when "101001010110" => A <= "000000000000000000"; -- Line 11   Column 87   Coefficient 0.00000000
         when "101001010111" => A <= "000000000000000000"; -- Line 11   Column 88   Coefficient 0.00000000
         when "101001011000" => A <= "000000000000000000"; -- Line 11   Column 89   Coefficient 0.00000000
         when "101001011001" => A <= "000000000000000000"; -- Line 11   Column 90   Coefficient 0.00000000
         when "101001011010" => A <= "000000000000000000"; -- Line 11   Column 91   Coefficient 0.00000000
         when "101001011011" => A <= "000000000000000000"; -- Line 11   Column 92   Coefficient 0.00000000
         when "101001011100" => A <= "000000000000000000"; -- Line 11   Column 93   Coefficient 0.00000000
         when "101001011101" => A <= "000000000000000000"; -- Line 11   Column 94   Coefficient 0.00000000
         when "101001011110" => A <= "000000000000000000"; -- Line 11   Column 95   Coefficient 0.00000000
         when "101001011111" => A <= "000000000000000000"; -- Line 11   Column 96   Coefficient 0.00000000
         when "101001100000" => A <= "000000000000000000"; -- Line 11   Column 97   Coefficient 0.00000000
         when "101001100001" => A <= "000000000000000000"; -- Line 11   Column 98   Coefficient 0.00000000
         when "101001100010" => A <= "000000000000000000"; -- Line 11   Column 99   Coefficient 0.00000000
         when "101001100011" => A <= "000000000000000000"; -- Line 11   Column 100   Coefficient 0.00000000
         when "101001100100" => A <= "000000000000000000"; -- Line 11   Column 101   Coefficient 0.00000000
         when "101001100101" => A <= "000000000000000000"; -- Line 11   Column 102   Coefficient 0.00000000
         when "101001100110" => A <= "000000000000000000"; -- Line 11   Column 103   Coefficient 0.00000000
         when "101001100111" => A <= "000000000000000000"; -- Line 11   Column 104   Coefficient 0.00000000
         when "101001101000" => A <= "000000000000000000"; -- Line 11   Column 105   Coefficient 0.00000000
         when "101001101001" => A <= "000000000000000000"; -- Line 11   Column 106   Coefficient 0.00000000
         when "101001101010" => A <= "000000000000000000"; -- Line 11   Column 107   Coefficient 0.00000000
         when "101001101011" => A <= "000000000000000000"; -- Line 11   Column 108   Coefficient 0.00000000
         when "101001101100" => A <= "000000000000000000"; -- Line 11   Column 109   Coefficient 0.00000000
         when "101001101101" => A <= "000000000000000000"; -- Line 11   Column 110   Coefficient 0.00000000
         when "101001101110" => A <= "000000000000000000"; -- Line 11   Column 111   Coefficient 0.00000000
         when "101001101111" => A <= "000000000000000000"; -- Line 11   Column 112   Coefficient 0.00000000
         when "101001110000" => A <= "000000000000000000"; -- Line 11   Column 113   Coefficient 0.00000000
         when "101001110001" => A <= "000000000000000000"; -- Line 11   Column 114   Coefficient 0.00000000
         when "101001110010" => A <= "000000000000000000"; -- Line 11   Column 115   Coefficient 0.00000000
         when "101001110011" => A <= "000000000000000000"; -- Line 11   Column 116   Coefficient 0.00000000
         when "101001110100" => A <= "000000000000000000"; -- Line 11   Column 117   Coefficient 0.00000000
         when "101001110101" => A <= "000000000000000000"; -- Line 11   Column 118   Coefficient 0.00000000
         when "101001110110" => A <= "000000000000000000"; -- Line 11   Column 119   Coefficient 0.00000000
         when "101001110111" => A <= "000000000000000000"; -- Line 11   Column 120   Coefficient 0.00000000
         when "101001111000" => A <= "000000000000000000"; -- Line 11   Column 121   Coefficient 0.00000000
         when "101001111001" => A <= "000000000000000000"; -- Line 11   Column 122   Coefficient 0.00000000
         when "101001111010" => A <= "000000000000000000"; -- Line 11   Column 123   Coefficient 0.00000000
         when "101001111011" => A <= "000000000000000000"; -- Line 11   Column 124   Coefficient 0.00000000
         when "101001111100" => A <= "000000000000000000"; -- Line 11   Column 125   Coefficient 0.00000000
         when "101001111101" => A <= "000000000000000000"; -- Line 11   Column 126   Coefficient 0.00000000
         when "101001111110" => A <= "000000000000000000"; -- Line 11   Column 127   Coefficient 0.00000000
         when "101001111111" => A <= "000000000000000000"; -- Line 11   Column 128   Coefficient 0.00000000
         when "101010000000" => A <= "000000000000000000"; -- Line 11   Column 129   Coefficient 0.00000000
         when "101010000001" => A <= "000000000000000000"; -- Line 11   Column 130   Coefficient 0.00000000
         when "101010000010" => A <= "000000000000000000"; -- Line 11   Column 131   Coefficient 0.00000000
         when "101010000011" => A <= "000000000000000000"; -- Line 11   Column 132   Coefficient 0.00000000
         when "101010000100" => A <= "000000000000000000"; -- Line 11   Column 133   Coefficient 0.00000000
         when "101010000101" => A <= "000000000000000000"; -- Line 11   Column 134   Coefficient 0.00000000
         when "101010000110" => A <= "000000000000000000"; -- Line 11   Column 135   Coefficient 0.00000000
         when "101010000111" => A <= "000000000000000000"; -- Line 11   Column 136   Coefficient 0.00000000
         when "101010001000" => A <= "000000000000000000"; -- Line 11   Column 137   Coefficient 0.00000000
         when "101010001001" => A <= "000000000000000000"; -- Line 11   Column 138   Coefficient 0.00000000
         when "101010001010" => A <= "000000000000000000"; -- Line 11   Column 139   Coefficient 0.00000000
         when "101010001011" => A <= "000000000000000000"; -- Line 11   Column 140   Coefficient 0.00000000
         when "101010001100" => A <= "000000000000000000"; -- Line 11   Column 141   Coefficient 0.00000000
         when "101010001101" => A <= "000000000000000000"; -- Line 11   Column 142   Coefficient 0.00000000
         when "101010001110" => A <= "000000000000000000"; -- Line 11   Column 143   Coefficient 0.00000000
         when "101010001111" => A <= "000000000000000000"; -- Line 11   Column 144   Coefficient 0.00000000
         when "101010010000" => A <= "000000000000000000"; -- Line 11   Column 145   Coefficient 0.00000000
         when "101010010001" => A <= "000000000000000000"; -- Line 11   Column 146   Coefficient 0.00000000
         when "101010010010" => A <= "000000000000000000"; -- Line 11   Column 147   Coefficient 0.00000000
         when "101010010011" => A <= "000000000000000000"; -- Line 11   Column 148   Coefficient 0.00000000
         when "101010010100" => A <= "000000000000000000"; -- Line 11   Column 149   Coefficient 0.00000000
         when "101010010101" => A <= "000000000000000000"; -- Line 11   Column 150   Coefficient 0.00000000
         when "101010010110" => A <= "000000000000000000"; -- Line 11   Column 151   Coefficient 0.00000000
         when "101010010111" => A <= "000000000000000000"; -- Line 11   Column 152   Coefficient 0.00000000
         when "101010011000" => A <= "000000000000000000"; -- Line 11   Column 153   Coefficient 0.00000000
         when "101010011001" => A <= "000000000000000000"; -- Line 11   Column 154   Coefficient 0.00000000
         when "101010011010" => A <= "000000000000000000"; -- Line 11   Column 155   Coefficient 0.00000000
         when "101010011011" => A <= "000000000000000000"; -- Line 11   Column 156   Coefficient 0.00000000
         when "101010011100" => A <= "000000000000000000"; -- Line 11   Column 157   Coefficient 0.00000000
         when "101010011101" => A <= "000000000000000000"; -- Line 11   Column 158   Coefficient 0.00000000
         when "101010011110" => A <= "000000000000000000"; -- Line 11   Column 159   Coefficient 0.00000000
         when "101010011111" => A <= "000000000000000000"; -- Line 11   Column 160   Coefficient 0.00000000
         when "101010100000" => A <= "000000000000001001"; -- Line 11   Column 161   Coefficient 0.00003433
         when "101010100001" => A <= "000000000000000011"; -- Line 11   Column 162   Coefficient 0.00001144
         when "101010100010" => A <= "111111111111001011"; -- Line 11   Column 163   Coefficient -0.00020218
         when "101010100011" => A <= "111111111110100110"; -- Line 11   Column 164   Coefficient -0.00034332
         when "101010100100" => A <= "111111111110010010"; -- Line 11   Column 165   Coefficient -0.00041962
         when "101010100101" => A <= "111111111111010011"; -- Line 11   Column 166   Coefficient -0.00017166
         when "101010100110" => A <= "000000000011111000"; -- Line 11   Column 167   Coefficient 0.00094604
         when "101010100111" => A <= "000000001000010011"; -- Line 11   Column 168   Coefficient 0.00202560
         when "101010101000" => A <= "000000001010110110"; -- Line 11   Column 169   Coefficient 0.00264740
         when "101010101001" => A <= "000000001101001100"; -- Line 11   Column 170   Coefficient 0.00321960
         when "101010101010" => A <= "000000001111111100"; -- Line 11   Column 171   Coefficient 0.00389099
         when "101010101011" => A <= "000000010000011000"; -- Line 11   Column 172   Coefficient 0.00399780
         when "101010101100" => A <= "000000001111000010"; -- Line 11   Column 173   Coefficient 0.00366974
         when "101010101101" => A <= "000000000111011010"; -- Line 11   Column 174   Coefficient 0.00180817
         when "101010101110" => A <= "111111110001010101"; -- Line 11   Column 175   Coefficient -0.00358200
         when "101010101111" => A <= "111111011001111001"; -- Line 11   Column 176   Coefficient -0.00930405
         when "101010110000" => A <= "111111000100111001"; -- Line 11   Column 177   Coefficient -0.01443100
         when "101010110001" => A <= "111110110001100001"; -- Line 11   Column 178   Coefficient -0.01916122
         when "101010110010" => A <= "111110100110010011"; -- Line 11   Column 179   Coefficient -0.02190018
         when "101010110011" => A <= "111110011011111010"; -- Line 11   Column 180   Coefficient -0.02443695
         when "101010110100" => A <= "111110010000110000"; -- Line 11   Column 181   Coefficient -0.02716064
         when "101010110101" => A <= "111110000101010011"; -- Line 11   Column 182   Coefficient -0.02995682
         when "101010110110" => A <= "111101110100001010"; -- Line 11   Column 183   Coefficient -0.03414154
         when "101010110111" => A <= "111101100110110000"; -- Line 11   Column 184   Coefficient -0.03741455
         when "101010111000" => A <= "111101100010101111"; -- Line 11   Column 185   Coefficient -0.03839493
         when "101010111001" => A <= "111101100010001110"; -- Line 11   Column 186   Coefficient -0.03852081
         when "101010111010" => A <= "111101100000101101"; -- Line 11   Column 187   Coefficient -0.03889084
         when "101010111011" => A <= "111101101011101110"; -- Line 11   Column 188   Coefficient -0.03620148
         when "101010111100" => A <= "111110000010011110"; -- Line 11   Column 189   Coefficient -0.03064728
         when "101010111101" => A <= "111110110101100100"; -- Line 11   Column 190   Coefficient -0.01817322
         when "101010111110" => A <= "000000100101011001"; -- Line 11   Column 191   Coefficient 0.00912857
         when "101010111111" => A <= "000010011110111100"; -- Line 11   Column 192   Coefficient 0.03880310
         when "101011000000" => A <= "000100010010000101"; -- Line 11   Column 193   Coefficient 0.06691360
         when "101011000001" => A <= "000110000101110011"; -- Line 11   Column 194   Coefficient 0.09516525
         when "101011000010" => A <= "000111100110110001"; -- Line 11   Column 195   Coefficient 0.11883926
         when "101011000011" => A <= "001001000110101001"; -- Line 11   Column 196   Coefficient 0.14224625
         when "101011000100" => A <= "001010101100000111"; -- Line 11   Column 197   Coefficient 0.16701889
         when "101011000101" => A <= "001100001011101000"; -- Line 11   Column 198   Coefficient 0.19033813
         when "101011000110" => A <= "001101100011111111"; -- Line 11   Column 199   Coefficient 0.21191025
         when "101011000111" => A <= "001110110101010100"; -- Line 11   Column 200   Coefficient 0.23176575
         when "101011001000" => A <= "001111111010100001"; -- Line 11   Column 201   Coefficient 0.24866104
         when "101011001001" => A <= "010000111010100101"; -- Line 11   Column 202   Coefficient 0.26430130
         when "101011001010" => A <= "010010000001100011"; -- Line 11   Column 203   Coefficient 0.28162766
         when "101011001011" => A <= "010010110100110100"; -- Line 11   Column 204   Coefficient 0.29414368
         when "101011001100" => A <= "010011010010100110"; -- Line 11   Column 205   Coefficient 0.30141449
         when "101011001101" => A <= "010011000101100111"; -- Line 11   Column 206   Coefficient 0.29824448
         when "101011001110" => A <= "010001011110001011"; -- Line 11   Column 207   Coefficient 0.27299118
         when "101011001111" => A <= "001111100101110011"; -- Line 11   Column 208   Coefficient 0.24360275
         when "101011010000" => A <= "001101110100101001"; -- Line 11   Column 209   Coefficient 0.21597672
         when "101011010001" => A <= "001011111101111010"; -- Line 11   Column 210   Coefficient 0.18698883
         when "101011010010" => A <= "001010011001111000"; -- Line 11   Column 211   Coefficient 0.16256714
         when "101011010011" => A <= "001000110101000000"; -- Line 11   Column 212   Coefficient 0.13793945
         when "101011010100" => A <= "000111000101010101"; -- Line 11   Column 213   Coefficient 0.11067581
         when "101011010101" => A <= "000101100000010101"; -- Line 11   Column 214   Coefficient 0.08601761
         when "101011010110" => A <= "000100010011001101"; -- Line 11   Column 215   Coefficient 0.06718826
         when "101011010111" => A <= "000011001010010011"; -- Line 11   Column 216   Coefficient 0.04938889
         when "101011011000" => A <= "000010000100001011"; -- Line 11   Column 217   Coefficient 0.03226852
         when "101011011001" => A <= "000000111110100110"; -- Line 11   Column 218   Coefficient 0.01528168
         when "101011011010" => A <= "111111101010001000"; -- Line 11   Column 219   Coefficient -0.00534058
         when "101011011011" => A <= "111110100000101100"; -- Line 11   Column 220   Coefficient -0.02326965
         when "101011011100" => A <= "111101100111001110"; -- Line 11   Column 221   Coefficient -0.03730011
         when "101011011101" => A <= "111101000110110001"; -- Line 11   Column 222   Coefficient -0.04522324
         when "101011011110" => A <= "111101011101101101"; -- Line 11   Column 223   Coefficient -0.03962326
         when "101011011111" => A <= "111101111110110001"; -- Line 11   Column 224   Coefficient -0.03155136
         when "101011100000" => A <= "111110011010010101"; -- Line 11   Column 225   Coefficient -0.02482224
         when "101011100001" => A <= "111110111010000001"; -- Line 11   Column 226   Coefficient -0.01708603
         when "101011100010" => A <= "111111010000101110"; -- Line 11   Column 227   Coefficient -0.01154327
         when "101011100011" => A <= "111111100111100010"; -- Line 11   Column 228   Coefficient -0.00597382
         when "101011100100" => A <= "000000000100100100"; -- Line 11   Column 229   Coefficient 0.00111389
         when "101011100101" => A <= "000000011000110111"; -- Line 11   Column 230   Coefficient 0.00606918
         when "101011100110" => A <= "000000010111101010"; -- Line 11   Column 231   Coefficient 0.00577545
         when "101011100111" => A <= "000000010100111001"; -- Line 11   Column 232   Coefficient 0.00510025
         when "101011101000" => A <= "000000010100110111"; -- Line 11   Column 233   Coefficient 0.00509262
         when "101011101001" => A <= "000000010110010000"; -- Line 11   Column 234   Coefficient 0.00543213
         when "101011101010" => A <= "000000100010100100"; -- Line 11   Column 235   Coefficient 0.00843811
         when "101011101011" => A <= "000000101101010111"; -- Line 11   Column 236   Coefficient 0.01107407
         when "101011101100" => A <= "000000110010101110"; -- Line 11   Column 237   Coefficient 0.01238251
         when "101011101101" => A <= "000000110100010110"; -- Line 11   Column 238   Coefficient 0.01277924
         when "101011101110" => A <= "000000101011110101"; -- Line 11   Column 239   Coefficient 0.01070023
         when "101011101111" => A <= "000000100001110011"; -- Line 11   Column 240   Coefficient 0.00825119
         when "101011110000" => A <= "000000011001110100"; -- Line 11   Column 241   Coefficient 0.00630188
         when "101011110001" => A <= "000000010001001000"; -- Line 11   Column 242   Coefficient 0.00418091
         when "101011110010" => A <= "000000001001011000"; -- Line 11   Column 243   Coefficient 0.00228882
         when "101011110011" => A <= "000000000010010011"; -- Line 11   Column 244   Coefficient 0.00056076
         when "101011110100" => A <= "111111111010111001"; -- Line 11   Column 245   Coefficient -0.00124741
         when "101011110101" => A <= "111111110110011111"; -- Line 11   Column 246   Coefficient -0.00232315
         when "101011110110" => A <= "111111111001000110"; -- Line 11   Column 247   Coefficient -0.00168610
         when "101011110111" => A <= "111111111100011110"; -- Line 11   Column 248   Coefficient -0.00086212
         when "101011111000" => A <= "111111111110110111"; -- Line 11   Column 249   Coefficient -0.00027847
         when "101011111001" => A <= "000000000001001011"; -- Line 11   Column 250   Coefficient 0.00028610
         when "101011111010" => A <= "000000000001001000"; -- Line 11   Column 251   Coefficient 0.00027466
         when "101011111011" => A <= "000000000001000010"; -- Line 11   Column 252   Coefficient 0.00025177
         when "101011111100" => A <= "000000000001111110"; -- Line 11   Column 253   Coefficient 0.00048065
         when "101011111101" => A <= "000000000010010101"; -- Line 11   Column 254   Coefficient 0.00056839
         when "101011111110" => A <= "000000000001100101"; -- Line 11   Column 255   Coefficient 0.00038528
         when "101011111111" => A <= "000000000000110011"; -- Line 11   Column 256   Coefficient 0.00019455
         when "101100000000" => A <= "000000011001110100"; -- Line 12   Column 1   Coefficient 0.00630188
         when "101100000001" => A <= "000000010001001000"; -- Line 12   Column 2   Coefficient 0.00418091
         when "101100000010" => A <= "000000001001011000"; -- Line 12   Column 3   Coefficient 0.00228882
         when "101100000011" => A <= "000000000010010011"; -- Line 12   Column 4   Coefficient 0.00056076
         when "101100000100" => A <= "111111111010111001"; -- Line 12   Column 5   Coefficient -0.00124741
         when "101100000101" => A <= "111111110110011111"; -- Line 12   Column 6   Coefficient -0.00232315
         when "101100000110" => A <= "111111111001000110"; -- Line 12   Column 7   Coefficient -0.00168610
         when "101100000111" => A <= "111111111100011110"; -- Line 12   Column 8   Coefficient -0.00086212
         when "101100001000" => A <= "111111111110110111"; -- Line 12   Column 9   Coefficient -0.00027847
         when "101100001001" => A <= "000000000001001011"; -- Line 12   Column 10   Coefficient 0.00028610
         when "101100001010" => A <= "000000000001001000"; -- Line 12   Column 11   Coefficient 0.00027466
         when "101100001011" => A <= "000000000001000010"; -- Line 12   Column 12   Coefficient 0.00025177
         when "101100001100" => A <= "000000000001111110"; -- Line 12   Column 13   Coefficient 0.00048065
         when "101100001101" => A <= "000000000010010101"; -- Line 12   Column 14   Coefficient 0.00056839
         when "101100001110" => A <= "000000000001100101"; -- Line 12   Column 15   Coefficient 0.00038528
         when "101100001111" => A <= "000000000000110011"; -- Line 12   Column 16   Coefficient 0.00019455
         when "101100010000" => A <= "000000000000000111"; -- Line 12   Column 17   Coefficient 0.00002670
         when "101100010001" => A <= "111111111111100110"; -- Line 12   Column 18   Coefficient -0.00009918
         when "101100010010" => A <= "111111111111110100"; -- Line 12   Column 19   Coefficient -0.00004578
         when "101100010011" => A <= "000000000000000011"; -- Line 12   Column 20   Coefficient 0.00001144
         when "101100010100" => A <= "000000000000000100"; -- Line 12   Column 21   Coefficient 0.00001526
         when "101100010101" => A <= "000000000000000110"; -- Line 12   Column 22   Coefficient 0.00002289
         when "101100010110" => A <= "000000000000000011"; -- Line 12   Column 23   Coefficient 0.00001144
         when "101100010111" => A <= "111111111111111111"; -- Line 12   Column 24   Coefficient -0.00000381
         when "101100011000" => A <= "000000000000000000"; -- Line 12   Column 25   Coefficient 0.00000000
         when "101100011001" => A <= "000000000000000000"; -- Line 12   Column 26   Coefficient 0.00000000
         when "101100011010" => A <= "000000000000000000"; -- Line 12   Column 27   Coefficient 0.00000000
         when "101100011011" => A <= "000000000000000000"; -- Line 12   Column 28   Coefficient 0.00000000
         when "101100011100" => A <= "000000000000000000"; -- Line 12   Column 29   Coefficient 0.00000000
         when "101100011101" => A <= "000000000000000000"; -- Line 12   Column 30   Coefficient 0.00000000
         when "101100011110" => A <= "000000000000000000"; -- Line 12   Column 31   Coefficient 0.00000000
         when "101100011111" => A <= "000000000000000000"; -- Line 12   Column 32   Coefficient 0.00000000
         when "101100100000" => A <= "000000000000000000"; -- Line 12   Column 33   Coefficient 0.00000000
         when "101100100001" => A <= "000000000000000000"; -- Line 12   Column 34   Coefficient 0.00000000
         when "101100100010" => A <= "000000000000000000"; -- Line 12   Column 35   Coefficient 0.00000000
         when "101100100011" => A <= "000000000000000000"; -- Line 12   Column 36   Coefficient 0.00000000
         when "101100100100" => A <= "000000000000000000"; -- Line 12   Column 37   Coefficient 0.00000000
         when "101100100101" => A <= "000000000000000000"; -- Line 12   Column 38   Coefficient 0.00000000
         when "101100100110" => A <= "000000000000000000"; -- Line 12   Column 39   Coefficient 0.00000000
         when "101100100111" => A <= "000000000000000000"; -- Line 12   Column 40   Coefficient 0.00000000
         when "101100101000" => A <= "000000000000000000"; -- Line 12   Column 41   Coefficient 0.00000000
         when "101100101001" => A <= "000000000000000000"; -- Line 12   Column 42   Coefficient 0.00000000
         when "101100101010" => A <= "000000000000000000"; -- Line 12   Column 43   Coefficient 0.00000000
         when "101100101011" => A <= "000000000000000000"; -- Line 12   Column 44   Coefficient 0.00000000
         when "101100101100" => A <= "000000000000000000"; -- Line 12   Column 45   Coefficient 0.00000000
         when "101100101101" => A <= "000000000000000000"; -- Line 12   Column 46   Coefficient 0.00000000
         when "101100101110" => A <= "000000000000000000"; -- Line 12   Column 47   Coefficient 0.00000000
         when "101100101111" => A <= "000000000000000000"; -- Line 12   Column 48   Coefficient 0.00000000
         when "101100110000" => A <= "000000000000000000"; -- Line 12   Column 49   Coefficient 0.00000000
         when "101100110001" => A <= "000000000000000000"; -- Line 12   Column 50   Coefficient 0.00000000
         when "101100110010" => A <= "000000000000000000"; -- Line 12   Column 51   Coefficient 0.00000000
         when "101100110011" => A <= "000000000000000000"; -- Line 12   Column 52   Coefficient 0.00000000
         when "101100110100" => A <= "000000000000000000"; -- Line 12   Column 53   Coefficient 0.00000000
         when "101100110101" => A <= "000000000000000000"; -- Line 12   Column 54   Coefficient 0.00000000
         when "101100110110" => A <= "000000000000000000"; -- Line 12   Column 55   Coefficient 0.00000000
         when "101100110111" => A <= "000000000000000000"; -- Line 12   Column 56   Coefficient 0.00000000
         when "101100111000" => A <= "000000000000000000"; -- Line 12   Column 57   Coefficient 0.00000000
         when "101100111001" => A <= "000000000000000000"; -- Line 12   Column 58   Coefficient 0.00000000
         when "101100111010" => A <= "000000000000000000"; -- Line 12   Column 59   Coefficient 0.00000000
         when "101100111011" => A <= "000000000000000000"; -- Line 12   Column 60   Coefficient 0.00000000
         when "101100111100" => A <= "000000000000000000"; -- Line 12   Column 61   Coefficient 0.00000000
         when "101100111101" => A <= "000000000000000000"; -- Line 12   Column 62   Coefficient 0.00000000
         when "101100111110" => A <= "000000000000000000"; -- Line 12   Column 63   Coefficient 0.00000000
         when "101100111111" => A <= "000000000000000000"; -- Line 12   Column 64   Coefficient 0.00000000
         when "101101000000" => A <= "000000000000000000"; -- Line 12   Column 65   Coefficient 0.00000000
         when "101101000001" => A <= "000000000000000000"; -- Line 12   Column 66   Coefficient 0.00000000
         when "101101000010" => A <= "000000000000000000"; -- Line 12   Column 67   Coefficient 0.00000000
         when "101101000011" => A <= "000000000000000000"; -- Line 12   Column 68   Coefficient 0.00000000
         when "101101000100" => A <= "000000000000000000"; -- Line 12   Column 69   Coefficient 0.00000000
         when "101101000101" => A <= "000000000000000000"; -- Line 12   Column 70   Coefficient 0.00000000
         when "101101000110" => A <= "000000000000000000"; -- Line 12   Column 71   Coefficient 0.00000000
         when "101101000111" => A <= "000000000000000000"; -- Line 12   Column 72   Coefficient 0.00000000
         when "101101001000" => A <= "000000000000000000"; -- Line 12   Column 73   Coefficient 0.00000000
         when "101101001001" => A <= "000000000000000000"; -- Line 12   Column 74   Coefficient 0.00000000
         when "101101001010" => A <= "000000000000000000"; -- Line 12   Column 75   Coefficient 0.00000000
         when "101101001011" => A <= "000000000000000000"; -- Line 12   Column 76   Coefficient 0.00000000
         when "101101001100" => A <= "000000000000000000"; -- Line 12   Column 77   Coefficient 0.00000000
         when "101101001101" => A <= "000000000000000000"; -- Line 12   Column 78   Coefficient 0.00000000
         when "101101001110" => A <= "000000000000000000"; -- Line 12   Column 79   Coefficient 0.00000000
         when "101101001111" => A <= "000000000000000000"; -- Line 12   Column 80   Coefficient 0.00000000
         when "101101010000" => A <= "000000000000000000"; -- Line 12   Column 81   Coefficient 0.00000000
         when "101101010001" => A <= "000000000000000000"; -- Line 12   Column 82   Coefficient 0.00000000
         when "101101010010" => A <= "000000000000000000"; -- Line 12   Column 83   Coefficient 0.00000000
         when "101101010011" => A <= "000000000000000000"; -- Line 12   Column 84   Coefficient 0.00000000
         when "101101010100" => A <= "000000000000000000"; -- Line 12   Column 85   Coefficient 0.00000000
         when "101101010101" => A <= "000000000000000000"; -- Line 12   Column 86   Coefficient 0.00000000
         when "101101010110" => A <= "000000000000000000"; -- Line 12   Column 87   Coefficient 0.00000000
         when "101101010111" => A <= "000000000000000000"; -- Line 12   Column 88   Coefficient 0.00000000
         when "101101011000" => A <= "000000000000000000"; -- Line 12   Column 89   Coefficient 0.00000000
         when "101101011001" => A <= "000000000000000000"; -- Line 12   Column 90   Coefficient 0.00000000
         when "101101011010" => A <= "000000000000000000"; -- Line 12   Column 91   Coefficient 0.00000000
         when "101101011011" => A <= "000000000000000000"; -- Line 12   Column 92   Coefficient 0.00000000
         when "101101011100" => A <= "000000000000000000"; -- Line 12   Column 93   Coefficient 0.00000000
         when "101101011101" => A <= "000000000000000000"; -- Line 12   Column 94   Coefficient 0.00000000
         when "101101011110" => A <= "000000000000000000"; -- Line 12   Column 95   Coefficient 0.00000000
         when "101101011111" => A <= "000000000000000000"; -- Line 12   Column 96   Coefficient 0.00000000
         when "101101100000" => A <= "000000000000000000"; -- Line 12   Column 97   Coefficient 0.00000000
         when "101101100001" => A <= "000000000000000000"; -- Line 12   Column 98   Coefficient 0.00000000
         when "101101100010" => A <= "000000000000000000"; -- Line 12   Column 99   Coefficient 0.00000000
         when "101101100011" => A <= "000000000000000000"; -- Line 12   Column 100   Coefficient 0.00000000
         when "101101100100" => A <= "000000000000000000"; -- Line 12   Column 101   Coefficient 0.00000000
         when "101101100101" => A <= "000000000000000000"; -- Line 12   Column 102   Coefficient 0.00000000
         when "101101100110" => A <= "000000000000000000"; -- Line 12   Column 103   Coefficient 0.00000000
         when "101101100111" => A <= "000000000000000000"; -- Line 12   Column 104   Coefficient 0.00000000
         when "101101101000" => A <= "000000000000000000"; -- Line 12   Column 105   Coefficient 0.00000000
         when "101101101001" => A <= "000000000000000000"; -- Line 12   Column 106   Coefficient 0.00000000
         when "101101101010" => A <= "000000000000000000"; -- Line 12   Column 107   Coefficient 0.00000000
         when "101101101011" => A <= "000000000000000000"; -- Line 12   Column 108   Coefficient 0.00000000
         when "101101101100" => A <= "000000000000000000"; -- Line 12   Column 109   Coefficient 0.00000000
         when "101101101101" => A <= "000000000000000000"; -- Line 12   Column 110   Coefficient 0.00000000
         when "101101101110" => A <= "000000000000000000"; -- Line 12   Column 111   Coefficient 0.00000000
         when "101101101111" => A <= "000000000000000000"; -- Line 12   Column 112   Coefficient 0.00000000
         when "101101110000" => A <= "000000000000000000"; -- Line 12   Column 113   Coefficient 0.00000000
         when "101101110001" => A <= "000000000000000000"; -- Line 12   Column 114   Coefficient 0.00000000
         when "101101110010" => A <= "000000000000000000"; -- Line 12   Column 115   Coefficient 0.00000000
         when "101101110011" => A <= "000000000000000000"; -- Line 12   Column 116   Coefficient 0.00000000
         when "101101110100" => A <= "000000000000000000"; -- Line 12   Column 117   Coefficient 0.00000000
         when "101101110101" => A <= "000000000000000000"; -- Line 12   Column 118   Coefficient 0.00000000
         when "101101110110" => A <= "000000000000000000"; -- Line 12   Column 119   Coefficient 0.00000000
         when "101101110111" => A <= "000000000000000000"; -- Line 12   Column 120   Coefficient 0.00000000
         when "101101111000" => A <= "000000000000000000"; -- Line 12   Column 121   Coefficient 0.00000000
         when "101101111001" => A <= "000000000000000000"; -- Line 12   Column 122   Coefficient 0.00000000
         when "101101111010" => A <= "000000000000000000"; -- Line 12   Column 123   Coefficient 0.00000000
         when "101101111011" => A <= "000000000000000000"; -- Line 12   Column 124   Coefficient 0.00000000
         when "101101111100" => A <= "000000000000000000"; -- Line 12   Column 125   Coefficient 0.00000000
         when "101101111101" => A <= "000000000000000000"; -- Line 12   Column 126   Coefficient 0.00000000
         when "101101111110" => A <= "000000000000000000"; -- Line 12   Column 127   Coefficient 0.00000000
         when "101101111111" => A <= "000000000000000000"; -- Line 12   Column 128   Coefficient 0.00000000
         when "101110000000" => A <= "000000000000000000"; -- Line 12   Column 129   Coefficient 0.00000000
         when "101110000001" => A <= "000000000000000000"; -- Line 12   Column 130   Coefficient 0.00000000
         when "101110000010" => A <= "000000000000000000"; -- Line 12   Column 131   Coefficient 0.00000000
         when "101110000011" => A <= "000000000000000000"; -- Line 12   Column 132   Coefficient 0.00000000
         when "101110000100" => A <= "000000000000000000"; -- Line 12   Column 133   Coefficient 0.00000000
         when "101110000101" => A <= "000000000000000000"; -- Line 12   Column 134   Coefficient 0.00000000
         when "101110000110" => A <= "000000000000000000"; -- Line 12   Column 135   Coefficient 0.00000000
         when "101110000111" => A <= "000000000000000000"; -- Line 12   Column 136   Coefficient 0.00000000
         when "101110001000" => A <= "000000000000000000"; -- Line 12   Column 137   Coefficient 0.00000000
         when "101110001001" => A <= "000000000000000000"; -- Line 12   Column 138   Coefficient 0.00000000
         when "101110001010" => A <= "000000000000000000"; -- Line 12   Column 139   Coefficient 0.00000000
         when "101110001011" => A <= "000000000000000000"; -- Line 12   Column 140   Coefficient 0.00000000
         when "101110001100" => A <= "000000000000000000"; -- Line 12   Column 141   Coefficient 0.00000000
         when "101110001101" => A <= "000000000000000000"; -- Line 12   Column 142   Coefficient 0.00000000
         when "101110001110" => A <= "000000000000000000"; -- Line 12   Column 143   Coefficient 0.00000000
         when "101110001111" => A <= "000000000000000000"; -- Line 12   Column 144   Coefficient 0.00000000
         when "101110010000" => A <= "000000000000000000"; -- Line 12   Column 145   Coefficient 0.00000000
         when "101110010001" => A <= "000000000000000000"; -- Line 12   Column 146   Coefficient 0.00000000
         when "101110010010" => A <= "000000000000000000"; -- Line 12   Column 147   Coefficient 0.00000000
         when "101110010011" => A <= "000000000000000000"; -- Line 12   Column 148   Coefficient 0.00000000
         when "101110010100" => A <= "000000000000000000"; -- Line 12   Column 149   Coefficient 0.00000000
         when "101110010101" => A <= "000000000000000000"; -- Line 12   Column 150   Coefficient 0.00000000
         when "101110010110" => A <= "000000000000000000"; -- Line 12   Column 151   Coefficient 0.00000000
         when "101110010111" => A <= "000000000000000000"; -- Line 12   Column 152   Coefficient 0.00000000
         when "101110011000" => A <= "000000000000000000"; -- Line 12   Column 153   Coefficient 0.00000000
         when "101110011001" => A <= "000000000000000000"; -- Line 12   Column 154   Coefficient 0.00000000
         when "101110011010" => A <= "000000000000000000"; -- Line 12   Column 155   Coefficient 0.00000000
         when "101110011011" => A <= "000000000000000000"; -- Line 12   Column 156   Coefficient 0.00000000
         when "101110011100" => A <= "000000000000000000"; -- Line 12   Column 157   Coefficient 0.00000000
         when "101110011101" => A <= "000000000000000000"; -- Line 12   Column 158   Coefficient 0.00000000
         when "101110011110" => A <= "000000000000000000"; -- Line 12   Column 159   Coefficient 0.00000000
         when "101110011111" => A <= "000000000000000000"; -- Line 12   Column 160   Coefficient 0.00000000
         when "101110100000" => A <= "000000000000000000"; -- Line 12   Column 161   Coefficient 0.00000000
         when "101110100001" => A <= "000000000000000000"; -- Line 12   Column 162   Coefficient 0.00000000
         when "101110100010" => A <= "000000000000000000"; -- Line 12   Column 163   Coefficient 0.00000000
         when "101110100011" => A <= "000000000000000000"; -- Line 12   Column 164   Coefficient 0.00000000
         when "101110100100" => A <= "000000000000000000"; -- Line 12   Column 165   Coefficient 0.00000000
         when "101110100101" => A <= "000000000000000000"; -- Line 12   Column 166   Coefficient 0.00000000
         when "101110100110" => A <= "000000000000000000"; -- Line 12   Column 167   Coefficient 0.00000000
         when "101110100111" => A <= "000000000000000000"; -- Line 12   Column 168   Coefficient 0.00000000
         when "101110101000" => A <= "000000000000000000"; -- Line 12   Column 169   Coefficient 0.00000000
         when "101110101001" => A <= "000000000000000000"; -- Line 12   Column 170   Coefficient 0.00000000
         when "101110101010" => A <= "000000000000000000"; -- Line 12   Column 171   Coefficient 0.00000000
         when "101110101011" => A <= "000000000000000000"; -- Line 12   Column 172   Coefficient 0.00000000
         when "101110101100" => A <= "000000000000000000"; -- Line 12   Column 173   Coefficient 0.00000000
         when "101110101101" => A <= "000000000000000000"; -- Line 12   Column 174   Coefficient 0.00000000
         when "101110101110" => A <= "000000000000000000"; -- Line 12   Column 175   Coefficient 0.00000000
         when "101110101111" => A <= "000000000000000000"; -- Line 12   Column 176   Coefficient 0.00000000
         when "101110110000" => A <= "000000000000001001"; -- Line 12   Column 177   Coefficient 0.00003433
         when "101110110001" => A <= "000000000000000011"; -- Line 12   Column 178   Coefficient 0.00001144
         when "101110110010" => A <= "111111111111001011"; -- Line 12   Column 179   Coefficient -0.00020218
         when "101110110011" => A <= "111111111110100110"; -- Line 12   Column 180   Coefficient -0.00034332
         when "101110110100" => A <= "111111111110010010"; -- Line 12   Column 181   Coefficient -0.00041962
         when "101110110101" => A <= "111111111111010011"; -- Line 12   Column 182   Coefficient -0.00017166
         when "101110110110" => A <= "000000000011111000"; -- Line 12   Column 183   Coefficient 0.00094604
         when "101110110111" => A <= "000000001000010011"; -- Line 12   Column 184   Coefficient 0.00202560
         when "101110111000" => A <= "000000001010110110"; -- Line 12   Column 185   Coefficient 0.00264740
         when "101110111001" => A <= "000000001101001100"; -- Line 12   Column 186   Coefficient 0.00321960
         when "101110111010" => A <= "000000001111111100"; -- Line 12   Column 187   Coefficient 0.00389099
         when "101110111011" => A <= "000000010000011000"; -- Line 12   Column 188   Coefficient 0.00399780
         when "101110111100" => A <= "000000001111000010"; -- Line 12   Column 189   Coefficient 0.00366974
         when "101110111101" => A <= "000000000111011010"; -- Line 12   Column 190   Coefficient 0.00180817
         when "101110111110" => A <= "111111110001010101"; -- Line 12   Column 191   Coefficient -0.00358200
         when "101110111111" => A <= "111111011001111001"; -- Line 12   Column 192   Coefficient -0.00930405
         when "101111000000" => A <= "111111000100111001"; -- Line 12   Column 193   Coefficient -0.01443100
         when "101111000001" => A <= "111110110001100001"; -- Line 12   Column 194   Coefficient -0.01916122
         when "101111000010" => A <= "111110100110010011"; -- Line 12   Column 195   Coefficient -0.02190018
         when "101111000011" => A <= "111110011011111010"; -- Line 12   Column 196   Coefficient -0.02443695
         when "101111000100" => A <= "111110010000110000"; -- Line 12   Column 197   Coefficient -0.02716064
         when "101111000101" => A <= "111110000101010011"; -- Line 12   Column 198   Coefficient -0.02995682
         when "101111000110" => A <= "111101110100001010"; -- Line 12   Column 199   Coefficient -0.03414154
         when "101111000111" => A <= "111101100110110000"; -- Line 12   Column 200   Coefficient -0.03741455
         when "101111001000" => A <= "111101100010101111"; -- Line 12   Column 201   Coefficient -0.03839493
         when "101111001001" => A <= "111101100010001110"; -- Line 12   Column 202   Coefficient -0.03852081
         when "101111001010" => A <= "111101100000101101"; -- Line 12   Column 203   Coefficient -0.03889084
         when "101111001011" => A <= "111101101011101110"; -- Line 12   Column 204   Coefficient -0.03620148
         when "101111001100" => A <= "111110000010011110"; -- Line 12   Column 205   Coefficient -0.03064728
         when "101111001101" => A <= "111110110101100100"; -- Line 12   Column 206   Coefficient -0.01817322
         when "101111001110" => A <= "000000100101011001"; -- Line 12   Column 207   Coefficient 0.00912857
         when "101111001111" => A <= "000010011110111100"; -- Line 12   Column 208   Coefficient 0.03880310
         when "101111010000" => A <= "000100010010000101"; -- Line 12   Column 209   Coefficient 0.06691360
         when "101111010001" => A <= "000110000101110011"; -- Line 12   Column 210   Coefficient 0.09516525
         when "101111010010" => A <= "000111100110110001"; -- Line 12   Column 211   Coefficient 0.11883926
         when "101111010011" => A <= "001001000110101001"; -- Line 12   Column 212   Coefficient 0.14224625
         when "101111010100" => A <= "001010101100000111"; -- Line 12   Column 213   Coefficient 0.16701889
         when "101111010101" => A <= "001100001011101000"; -- Line 12   Column 214   Coefficient 0.19033813
         when "101111010110" => A <= "001101100011111111"; -- Line 12   Column 215   Coefficient 0.21191025
         when "101111010111" => A <= "001110110101010100"; -- Line 12   Column 216   Coefficient 0.23176575
         when "101111011000" => A <= "001111111010100001"; -- Line 12   Column 217   Coefficient 0.24866104
         when "101111011001" => A <= "010000111010100101"; -- Line 12   Column 218   Coefficient 0.26430130
         when "101111011010" => A <= "010010000001100011"; -- Line 12   Column 219   Coefficient 0.28162766
         when "101111011011" => A <= "010010110100110100"; -- Line 12   Column 220   Coefficient 0.29414368
         when "101111011100" => A <= "010011010010100110"; -- Line 12   Column 221   Coefficient 0.30141449
         when "101111011101" => A <= "010011000101100111"; -- Line 12   Column 222   Coefficient 0.29824448
         when "101111011110" => A <= "010001011110001011"; -- Line 12   Column 223   Coefficient 0.27299118
         when "101111011111" => A <= "001111100101110011"; -- Line 12   Column 224   Coefficient 0.24360275
         when "101111100000" => A <= "001101110100101001"; -- Line 12   Column 225   Coefficient 0.21597672
         when "101111100001" => A <= "001011111101111010"; -- Line 12   Column 226   Coefficient 0.18698883
         when "101111100010" => A <= "001010011001111000"; -- Line 12   Column 227   Coefficient 0.16256714
         when "101111100011" => A <= "001000110101000000"; -- Line 12   Column 228   Coefficient 0.13793945
         when "101111100100" => A <= "000111000101010101"; -- Line 12   Column 229   Coefficient 0.11067581
         when "101111100101" => A <= "000101100000010101"; -- Line 12   Column 230   Coefficient 0.08601761
         when "101111100110" => A <= "000100010011001101"; -- Line 12   Column 231   Coefficient 0.06718826
         when "101111100111" => A <= "000011001010010011"; -- Line 12   Column 232   Coefficient 0.04938889
         when "101111101000" => A <= "000010000100001011"; -- Line 12   Column 233   Coefficient 0.03226852
         when "101111101001" => A <= "000000111110100110"; -- Line 12   Column 234   Coefficient 0.01528168
         when "101111101010" => A <= "111111101010001000"; -- Line 12   Column 235   Coefficient -0.00534058
         when "101111101011" => A <= "111110100000101100"; -- Line 12   Column 236   Coefficient -0.02326965
         when "101111101100" => A <= "111101100111001110"; -- Line 12   Column 237   Coefficient -0.03730011
         when "101111101101" => A <= "111101000110110001"; -- Line 12   Column 238   Coefficient -0.04522324
         when "101111101110" => A <= "111101011101101101"; -- Line 12   Column 239   Coefficient -0.03962326
         when "101111101111" => A <= "111101111110110001"; -- Line 12   Column 240   Coefficient -0.03155136
         when "101111110000" => A <= "111110011010010101"; -- Line 12   Column 241   Coefficient -0.02482224
         when "101111110001" => A <= "111110111010000001"; -- Line 12   Column 242   Coefficient -0.01708603
         when "101111110010" => A <= "111111010000101110"; -- Line 12   Column 243   Coefficient -0.01154327
         when "101111110011" => A <= "111111100111100010"; -- Line 12   Column 244   Coefficient -0.00597382
         when "101111110100" => A <= "000000000100100100"; -- Line 12   Column 245   Coefficient 0.00111389
         when "101111110101" => A <= "000000011000110111"; -- Line 12   Column 246   Coefficient 0.00606918
         when "101111110110" => A <= "000000010111101010"; -- Line 12   Column 247   Coefficient 0.00577545
         when "101111110111" => A <= "000000010100111001"; -- Line 12   Column 248   Coefficient 0.00510025
         when "101111111000" => A <= "000000010100110111"; -- Line 12   Column 249   Coefficient 0.00509262
         when "101111111001" => A <= "000000010110010000"; -- Line 12   Column 250   Coefficient 0.00543213
         when "101111111010" => A <= "000000100010100100"; -- Line 12   Column 251   Coefficient 0.00843811
         when "101111111011" => A <= "000000101101010111"; -- Line 12   Column 252   Coefficient 0.01107407
         when "101111111100" => A <= "000000110010101110"; -- Line 12   Column 253   Coefficient 0.01238251
         when "101111111101" => A <= "000000110100010110"; -- Line 12   Column 254   Coefficient 0.01277924
         when "101111111110" => A <= "000000101011110101"; -- Line 12   Column 255   Coefficient 0.01070023
         when "101111111111" => A <= "000000100001110011"; -- Line 12   Column 256   Coefficient 0.00825119
         when "110000000000" => A <= "111110011010010101"; -- Line 13   Column 1   Coefficient -0.02482224
         when "110000000001" => A <= "111110111010000001"; -- Line 13   Column 2   Coefficient -0.01708603
         when "110000000010" => A <= "111111010000101110"; -- Line 13   Column 3   Coefficient -0.01154327
         when "110000000011" => A <= "111111100111100010"; -- Line 13   Column 4   Coefficient -0.00597382
         when "110000000100" => A <= "000000000100100100"; -- Line 13   Column 5   Coefficient 0.00111389
         when "110000000101" => A <= "000000011000110111"; -- Line 13   Column 6   Coefficient 0.00606918
         when "110000000110" => A <= "000000010111101010"; -- Line 13   Column 7   Coefficient 0.00577545
         when "110000000111" => A <= "000000010100111001"; -- Line 13   Column 8   Coefficient 0.00510025
         when "110000001000" => A <= "000000010100110111"; -- Line 13   Column 9   Coefficient 0.00509262
         when "110000001001" => A <= "000000010110010000"; -- Line 13   Column 10   Coefficient 0.00543213
         when "110000001010" => A <= "000000100010100100"; -- Line 13   Column 11   Coefficient 0.00843811
         when "110000001011" => A <= "000000101101010111"; -- Line 13   Column 12   Coefficient 0.01107407
         when "110000001100" => A <= "000000110010101110"; -- Line 13   Column 13   Coefficient 0.01238251
         when "110000001101" => A <= "000000110100010110"; -- Line 13   Column 14   Coefficient 0.01277924
         when "110000001110" => A <= "000000101011110101"; -- Line 13   Column 15   Coefficient 0.01070023
         when "110000001111" => A <= "000000100001110011"; -- Line 13   Column 16   Coefficient 0.00825119
         when "110000010000" => A <= "000000011001110100"; -- Line 13   Column 17   Coefficient 0.00630188
         when "110000010001" => A <= "000000010001001000"; -- Line 13   Column 18   Coefficient 0.00418091
         when "110000010010" => A <= "000000001001011000"; -- Line 13   Column 19   Coefficient 0.00228882
         when "110000010011" => A <= "000000000010010011"; -- Line 13   Column 20   Coefficient 0.00056076
         when "110000010100" => A <= "111111111010111001"; -- Line 13   Column 21   Coefficient -0.00124741
         when "110000010101" => A <= "111111110110011111"; -- Line 13   Column 22   Coefficient -0.00232315
         when "110000010110" => A <= "111111111001000110"; -- Line 13   Column 23   Coefficient -0.00168610
         when "110000010111" => A <= "111111111100011110"; -- Line 13   Column 24   Coefficient -0.00086212
         when "110000011000" => A <= "111111111110110111"; -- Line 13   Column 25   Coefficient -0.00027847
         when "110000011001" => A <= "000000000001001011"; -- Line 13   Column 26   Coefficient 0.00028610
         when "110000011010" => A <= "000000000001001000"; -- Line 13   Column 27   Coefficient 0.00027466
         when "110000011011" => A <= "000000000001000010"; -- Line 13   Column 28   Coefficient 0.00025177
         when "110000011100" => A <= "000000000001111110"; -- Line 13   Column 29   Coefficient 0.00048065
         when "110000011101" => A <= "000000000010010101"; -- Line 13   Column 30   Coefficient 0.00056839
         when "110000011110" => A <= "000000000001100101"; -- Line 13   Column 31   Coefficient 0.00038528
         when "110000011111" => A <= "000000000000110011"; -- Line 13   Column 32   Coefficient 0.00019455
         when "110000100000" => A <= "000000000000000111"; -- Line 13   Column 33   Coefficient 0.00002670
         when "110000100001" => A <= "111111111111100110"; -- Line 13   Column 34   Coefficient -0.00009918
         when "110000100010" => A <= "111111111111110100"; -- Line 13   Column 35   Coefficient -0.00004578
         when "110000100011" => A <= "000000000000000011"; -- Line 13   Column 36   Coefficient 0.00001144
         when "110000100100" => A <= "000000000000000100"; -- Line 13   Column 37   Coefficient 0.00001526
         when "110000100101" => A <= "000000000000000110"; -- Line 13   Column 38   Coefficient 0.00002289
         when "110000100110" => A <= "000000000000000011"; -- Line 13   Column 39   Coefficient 0.00001144
         when "110000100111" => A <= "111111111111111111"; -- Line 13   Column 40   Coefficient -0.00000381
         when "110000101000" => A <= "000000000000000000"; -- Line 13   Column 41   Coefficient 0.00000000
         when "110000101001" => A <= "000000000000000000"; -- Line 13   Column 42   Coefficient 0.00000000
         when "110000101010" => A <= "000000000000000000"; -- Line 13   Column 43   Coefficient 0.00000000
         when "110000101011" => A <= "000000000000000000"; -- Line 13   Column 44   Coefficient 0.00000000
         when "110000101100" => A <= "000000000000000000"; -- Line 13   Column 45   Coefficient 0.00000000
         when "110000101101" => A <= "000000000000000000"; -- Line 13   Column 46   Coefficient 0.00000000
         when "110000101110" => A <= "000000000000000000"; -- Line 13   Column 47   Coefficient 0.00000000
         when "110000101111" => A <= "000000000000000000"; -- Line 13   Column 48   Coefficient 0.00000000
         when "110000110000" => A <= "000000000000000000"; -- Line 13   Column 49   Coefficient 0.00000000
         when "110000110001" => A <= "000000000000000000"; -- Line 13   Column 50   Coefficient 0.00000000
         when "110000110010" => A <= "000000000000000000"; -- Line 13   Column 51   Coefficient 0.00000000
         when "110000110011" => A <= "000000000000000000"; -- Line 13   Column 52   Coefficient 0.00000000
         when "110000110100" => A <= "000000000000000000"; -- Line 13   Column 53   Coefficient 0.00000000
         when "110000110101" => A <= "000000000000000000"; -- Line 13   Column 54   Coefficient 0.00000000
         when "110000110110" => A <= "000000000000000000"; -- Line 13   Column 55   Coefficient 0.00000000
         when "110000110111" => A <= "000000000000000000"; -- Line 13   Column 56   Coefficient 0.00000000
         when "110000111000" => A <= "000000000000000000"; -- Line 13   Column 57   Coefficient 0.00000000
         when "110000111001" => A <= "000000000000000000"; -- Line 13   Column 58   Coefficient 0.00000000
         when "110000111010" => A <= "000000000000000000"; -- Line 13   Column 59   Coefficient 0.00000000
         when "110000111011" => A <= "000000000000000000"; -- Line 13   Column 60   Coefficient 0.00000000
         when "110000111100" => A <= "000000000000000000"; -- Line 13   Column 61   Coefficient 0.00000000
         when "110000111101" => A <= "000000000000000000"; -- Line 13   Column 62   Coefficient 0.00000000
         when "110000111110" => A <= "000000000000000000"; -- Line 13   Column 63   Coefficient 0.00000000
         when "110000111111" => A <= "000000000000000000"; -- Line 13   Column 64   Coefficient 0.00000000
         when "110001000000" => A <= "000000000000000000"; -- Line 13   Column 65   Coefficient 0.00000000
         when "110001000001" => A <= "000000000000000000"; -- Line 13   Column 66   Coefficient 0.00000000
         when "110001000010" => A <= "000000000000000000"; -- Line 13   Column 67   Coefficient 0.00000000
         when "110001000011" => A <= "000000000000000000"; -- Line 13   Column 68   Coefficient 0.00000000
         when "110001000100" => A <= "000000000000000000"; -- Line 13   Column 69   Coefficient 0.00000000
         when "110001000101" => A <= "000000000000000000"; -- Line 13   Column 70   Coefficient 0.00000000
         when "110001000110" => A <= "000000000000000000"; -- Line 13   Column 71   Coefficient 0.00000000
         when "110001000111" => A <= "000000000000000000"; -- Line 13   Column 72   Coefficient 0.00000000
         when "110001001000" => A <= "000000000000000000"; -- Line 13   Column 73   Coefficient 0.00000000
         when "110001001001" => A <= "000000000000000000"; -- Line 13   Column 74   Coefficient 0.00000000
         when "110001001010" => A <= "000000000000000000"; -- Line 13   Column 75   Coefficient 0.00000000
         when "110001001011" => A <= "000000000000000000"; -- Line 13   Column 76   Coefficient 0.00000000
         when "110001001100" => A <= "000000000000000000"; -- Line 13   Column 77   Coefficient 0.00000000
         when "110001001101" => A <= "000000000000000000"; -- Line 13   Column 78   Coefficient 0.00000000
         when "110001001110" => A <= "000000000000000000"; -- Line 13   Column 79   Coefficient 0.00000000
         when "110001001111" => A <= "000000000000000000"; -- Line 13   Column 80   Coefficient 0.00000000
         when "110001010000" => A <= "000000000000000000"; -- Line 13   Column 81   Coefficient 0.00000000
         when "110001010001" => A <= "000000000000000000"; -- Line 13   Column 82   Coefficient 0.00000000
         when "110001010010" => A <= "000000000000000000"; -- Line 13   Column 83   Coefficient 0.00000000
         when "110001010011" => A <= "000000000000000000"; -- Line 13   Column 84   Coefficient 0.00000000
         when "110001010100" => A <= "000000000000000000"; -- Line 13   Column 85   Coefficient 0.00000000
         when "110001010101" => A <= "000000000000000000"; -- Line 13   Column 86   Coefficient 0.00000000
         when "110001010110" => A <= "000000000000000000"; -- Line 13   Column 87   Coefficient 0.00000000
         when "110001010111" => A <= "000000000000000000"; -- Line 13   Column 88   Coefficient 0.00000000
         when "110001011000" => A <= "000000000000000000"; -- Line 13   Column 89   Coefficient 0.00000000
         when "110001011001" => A <= "000000000000000000"; -- Line 13   Column 90   Coefficient 0.00000000
         when "110001011010" => A <= "000000000000000000"; -- Line 13   Column 91   Coefficient 0.00000000
         when "110001011011" => A <= "000000000000000000"; -- Line 13   Column 92   Coefficient 0.00000000
         when "110001011100" => A <= "000000000000000000"; -- Line 13   Column 93   Coefficient 0.00000000
         when "110001011101" => A <= "000000000000000000"; -- Line 13   Column 94   Coefficient 0.00000000
         when "110001011110" => A <= "000000000000000000"; -- Line 13   Column 95   Coefficient 0.00000000
         when "110001011111" => A <= "000000000000000000"; -- Line 13   Column 96   Coefficient 0.00000000
         when "110001100000" => A <= "000000000000000000"; -- Line 13   Column 97   Coefficient 0.00000000
         when "110001100001" => A <= "000000000000000000"; -- Line 13   Column 98   Coefficient 0.00000000
         when "110001100010" => A <= "000000000000000000"; -- Line 13   Column 99   Coefficient 0.00000000
         when "110001100011" => A <= "000000000000000000"; -- Line 13   Column 100   Coefficient 0.00000000
         when "110001100100" => A <= "000000000000000000"; -- Line 13   Column 101   Coefficient 0.00000000
         when "110001100101" => A <= "000000000000000000"; -- Line 13   Column 102   Coefficient 0.00000000
         when "110001100110" => A <= "000000000000000000"; -- Line 13   Column 103   Coefficient 0.00000000
         when "110001100111" => A <= "000000000000000000"; -- Line 13   Column 104   Coefficient 0.00000000
         when "110001101000" => A <= "000000000000000000"; -- Line 13   Column 105   Coefficient 0.00000000
         when "110001101001" => A <= "000000000000000000"; -- Line 13   Column 106   Coefficient 0.00000000
         when "110001101010" => A <= "000000000000000000"; -- Line 13   Column 107   Coefficient 0.00000000
         when "110001101011" => A <= "000000000000000000"; -- Line 13   Column 108   Coefficient 0.00000000
         when "110001101100" => A <= "000000000000000000"; -- Line 13   Column 109   Coefficient 0.00000000
         when "110001101101" => A <= "000000000000000000"; -- Line 13   Column 110   Coefficient 0.00000000
         when "110001101110" => A <= "000000000000000000"; -- Line 13   Column 111   Coefficient 0.00000000
         when "110001101111" => A <= "000000000000000000"; -- Line 13   Column 112   Coefficient 0.00000000
         when "110001110000" => A <= "000000000000000000"; -- Line 13   Column 113   Coefficient 0.00000000
         when "110001110001" => A <= "000000000000000000"; -- Line 13   Column 114   Coefficient 0.00000000
         when "110001110010" => A <= "000000000000000000"; -- Line 13   Column 115   Coefficient 0.00000000
         when "110001110011" => A <= "000000000000000000"; -- Line 13   Column 116   Coefficient 0.00000000
         when "110001110100" => A <= "000000000000000000"; -- Line 13   Column 117   Coefficient 0.00000000
         when "110001110101" => A <= "000000000000000000"; -- Line 13   Column 118   Coefficient 0.00000000
         when "110001110110" => A <= "000000000000000000"; -- Line 13   Column 119   Coefficient 0.00000000
         when "110001110111" => A <= "000000000000000000"; -- Line 13   Column 120   Coefficient 0.00000000
         when "110001111000" => A <= "000000000000000000"; -- Line 13   Column 121   Coefficient 0.00000000
         when "110001111001" => A <= "000000000000000000"; -- Line 13   Column 122   Coefficient 0.00000000
         when "110001111010" => A <= "000000000000000000"; -- Line 13   Column 123   Coefficient 0.00000000
         when "110001111011" => A <= "000000000000000000"; -- Line 13   Column 124   Coefficient 0.00000000
         when "110001111100" => A <= "000000000000000000"; -- Line 13   Column 125   Coefficient 0.00000000
         when "110001111101" => A <= "000000000000000000"; -- Line 13   Column 126   Coefficient 0.00000000
         when "110001111110" => A <= "000000000000000000"; -- Line 13   Column 127   Coefficient 0.00000000
         when "110001111111" => A <= "000000000000000000"; -- Line 13   Column 128   Coefficient 0.00000000
         when "110010000000" => A <= "000000000000000000"; -- Line 13   Column 129   Coefficient 0.00000000
         when "110010000001" => A <= "000000000000000000"; -- Line 13   Column 130   Coefficient 0.00000000
         when "110010000010" => A <= "000000000000000000"; -- Line 13   Column 131   Coefficient 0.00000000
         when "110010000011" => A <= "000000000000000000"; -- Line 13   Column 132   Coefficient 0.00000000
         when "110010000100" => A <= "000000000000000000"; -- Line 13   Column 133   Coefficient 0.00000000
         when "110010000101" => A <= "000000000000000000"; -- Line 13   Column 134   Coefficient 0.00000000
         when "110010000110" => A <= "000000000000000000"; -- Line 13   Column 135   Coefficient 0.00000000
         when "110010000111" => A <= "000000000000000000"; -- Line 13   Column 136   Coefficient 0.00000000
         when "110010001000" => A <= "000000000000000000"; -- Line 13   Column 137   Coefficient 0.00000000
         when "110010001001" => A <= "000000000000000000"; -- Line 13   Column 138   Coefficient 0.00000000
         when "110010001010" => A <= "000000000000000000"; -- Line 13   Column 139   Coefficient 0.00000000
         when "110010001011" => A <= "000000000000000000"; -- Line 13   Column 140   Coefficient 0.00000000
         when "110010001100" => A <= "000000000000000000"; -- Line 13   Column 141   Coefficient 0.00000000
         when "110010001101" => A <= "000000000000000000"; -- Line 13   Column 142   Coefficient 0.00000000
         when "110010001110" => A <= "000000000000000000"; -- Line 13   Column 143   Coefficient 0.00000000
         when "110010001111" => A <= "000000000000000000"; -- Line 13   Column 144   Coefficient 0.00000000
         when "110010010000" => A <= "000000000000000000"; -- Line 13   Column 145   Coefficient 0.00000000
         when "110010010001" => A <= "000000000000000000"; -- Line 13   Column 146   Coefficient 0.00000000
         when "110010010010" => A <= "000000000000000000"; -- Line 13   Column 147   Coefficient 0.00000000
         when "110010010011" => A <= "000000000000000000"; -- Line 13   Column 148   Coefficient 0.00000000
         when "110010010100" => A <= "000000000000000000"; -- Line 13   Column 149   Coefficient 0.00000000
         when "110010010101" => A <= "000000000000000000"; -- Line 13   Column 150   Coefficient 0.00000000
         when "110010010110" => A <= "000000000000000000"; -- Line 13   Column 151   Coefficient 0.00000000
         when "110010010111" => A <= "000000000000000000"; -- Line 13   Column 152   Coefficient 0.00000000
         when "110010011000" => A <= "000000000000000000"; -- Line 13   Column 153   Coefficient 0.00000000
         when "110010011001" => A <= "000000000000000000"; -- Line 13   Column 154   Coefficient 0.00000000
         when "110010011010" => A <= "000000000000000000"; -- Line 13   Column 155   Coefficient 0.00000000
         when "110010011011" => A <= "000000000000000000"; -- Line 13   Column 156   Coefficient 0.00000000
         when "110010011100" => A <= "000000000000000000"; -- Line 13   Column 157   Coefficient 0.00000000
         when "110010011101" => A <= "000000000000000000"; -- Line 13   Column 158   Coefficient 0.00000000
         when "110010011110" => A <= "000000000000000000"; -- Line 13   Column 159   Coefficient 0.00000000
         when "110010011111" => A <= "000000000000000000"; -- Line 13   Column 160   Coefficient 0.00000000
         when "110010100000" => A <= "000000000000000000"; -- Line 13   Column 161   Coefficient 0.00000000
         when "110010100001" => A <= "000000000000000000"; -- Line 13   Column 162   Coefficient 0.00000000
         when "110010100010" => A <= "000000000000000000"; -- Line 13   Column 163   Coefficient 0.00000000
         when "110010100011" => A <= "000000000000000000"; -- Line 13   Column 164   Coefficient 0.00000000
         when "110010100100" => A <= "000000000000000000"; -- Line 13   Column 165   Coefficient 0.00000000
         when "110010100101" => A <= "000000000000000000"; -- Line 13   Column 166   Coefficient 0.00000000
         when "110010100110" => A <= "000000000000000000"; -- Line 13   Column 167   Coefficient 0.00000000
         when "110010100111" => A <= "000000000000000000"; -- Line 13   Column 168   Coefficient 0.00000000
         when "110010101000" => A <= "000000000000000000"; -- Line 13   Column 169   Coefficient 0.00000000
         when "110010101001" => A <= "000000000000000000"; -- Line 13   Column 170   Coefficient 0.00000000
         when "110010101010" => A <= "000000000000000000"; -- Line 13   Column 171   Coefficient 0.00000000
         when "110010101011" => A <= "000000000000000000"; -- Line 13   Column 172   Coefficient 0.00000000
         when "110010101100" => A <= "000000000000000000"; -- Line 13   Column 173   Coefficient 0.00000000
         when "110010101101" => A <= "000000000000000000"; -- Line 13   Column 174   Coefficient 0.00000000
         when "110010101110" => A <= "000000000000000000"; -- Line 13   Column 175   Coefficient 0.00000000
         when "110010101111" => A <= "000000000000000000"; -- Line 13   Column 176   Coefficient 0.00000000
         when "110010110000" => A <= "000000000000000000"; -- Line 13   Column 177   Coefficient 0.00000000
         when "110010110001" => A <= "000000000000000000"; -- Line 13   Column 178   Coefficient 0.00000000
         when "110010110010" => A <= "000000000000000000"; -- Line 13   Column 179   Coefficient 0.00000000
         when "110010110011" => A <= "000000000000000000"; -- Line 13   Column 180   Coefficient 0.00000000
         when "110010110100" => A <= "000000000000000000"; -- Line 13   Column 181   Coefficient 0.00000000
         when "110010110101" => A <= "000000000000000000"; -- Line 13   Column 182   Coefficient 0.00000000
         when "110010110110" => A <= "000000000000000000"; -- Line 13   Column 183   Coefficient 0.00000000
         when "110010110111" => A <= "000000000000000000"; -- Line 13   Column 184   Coefficient 0.00000000
         when "110010111000" => A <= "000000000000000000"; -- Line 13   Column 185   Coefficient 0.00000000
         when "110010111001" => A <= "000000000000000000"; -- Line 13   Column 186   Coefficient 0.00000000
         when "110010111010" => A <= "000000000000000000"; -- Line 13   Column 187   Coefficient 0.00000000
         when "110010111011" => A <= "000000000000000000"; -- Line 13   Column 188   Coefficient 0.00000000
         when "110010111100" => A <= "000000000000000000"; -- Line 13   Column 189   Coefficient 0.00000000
         when "110010111101" => A <= "000000000000000000"; -- Line 13   Column 190   Coefficient 0.00000000
         when "110010111110" => A <= "000000000000000000"; -- Line 13   Column 191   Coefficient 0.00000000
         when "110010111111" => A <= "000000000000000000"; -- Line 13   Column 192   Coefficient 0.00000000
         when "110011000000" => A <= "000000000000001001"; -- Line 13   Column 193   Coefficient 0.00003433
         when "110011000001" => A <= "000000000000000011"; -- Line 13   Column 194   Coefficient 0.00001144
         when "110011000010" => A <= "111111111111001011"; -- Line 13   Column 195   Coefficient -0.00020218
         when "110011000011" => A <= "111111111110100110"; -- Line 13   Column 196   Coefficient -0.00034332
         when "110011000100" => A <= "111111111110010010"; -- Line 13   Column 197   Coefficient -0.00041962
         when "110011000101" => A <= "111111111111010011"; -- Line 13   Column 198   Coefficient -0.00017166
         when "110011000110" => A <= "000000000011111000"; -- Line 13   Column 199   Coefficient 0.00094604
         when "110011000111" => A <= "000000001000010011"; -- Line 13   Column 200   Coefficient 0.00202560
         when "110011001000" => A <= "000000001010110110"; -- Line 13   Column 201   Coefficient 0.00264740
         when "110011001001" => A <= "000000001101001100"; -- Line 13   Column 202   Coefficient 0.00321960
         when "110011001010" => A <= "000000001111111100"; -- Line 13   Column 203   Coefficient 0.00389099
         when "110011001011" => A <= "000000010000011000"; -- Line 13   Column 204   Coefficient 0.00399780
         when "110011001100" => A <= "000000001111000010"; -- Line 13   Column 205   Coefficient 0.00366974
         when "110011001101" => A <= "000000000111011010"; -- Line 13   Column 206   Coefficient 0.00180817
         when "110011001110" => A <= "111111110001010101"; -- Line 13   Column 207   Coefficient -0.00358200
         when "110011001111" => A <= "111111011001111001"; -- Line 13   Column 208   Coefficient -0.00930405
         when "110011010000" => A <= "111111000100111001"; -- Line 13   Column 209   Coefficient -0.01443100
         when "110011010001" => A <= "111110110001100001"; -- Line 13   Column 210   Coefficient -0.01916122
         when "110011010010" => A <= "111110100110010011"; -- Line 13   Column 211   Coefficient -0.02190018
         when "110011010011" => A <= "111110011011111010"; -- Line 13   Column 212   Coefficient -0.02443695
         when "110011010100" => A <= "111110010000110000"; -- Line 13   Column 213   Coefficient -0.02716064
         when "110011010101" => A <= "111110000101010011"; -- Line 13   Column 214   Coefficient -0.02995682
         when "110011010110" => A <= "111101110100001010"; -- Line 13   Column 215   Coefficient -0.03414154
         when "110011010111" => A <= "111101100110110000"; -- Line 13   Column 216   Coefficient -0.03741455
         when "110011011000" => A <= "111101100010101111"; -- Line 13   Column 217   Coefficient -0.03839493
         when "110011011001" => A <= "111101100010001110"; -- Line 13   Column 218   Coefficient -0.03852081
         when "110011011010" => A <= "111101100000101101"; -- Line 13   Column 219   Coefficient -0.03889084
         when "110011011011" => A <= "111101101011101110"; -- Line 13   Column 220   Coefficient -0.03620148
         when "110011011100" => A <= "111110000010011110"; -- Line 13   Column 221   Coefficient -0.03064728
         when "110011011101" => A <= "111110110101100100"; -- Line 13   Column 222   Coefficient -0.01817322
         when "110011011110" => A <= "000000100101011001"; -- Line 13   Column 223   Coefficient 0.00912857
         when "110011011111" => A <= "000010011110111100"; -- Line 13   Column 224   Coefficient 0.03880310
         when "110011100000" => A <= "000100010010000101"; -- Line 13   Column 225   Coefficient 0.06691360
         when "110011100001" => A <= "000110000101110011"; -- Line 13   Column 226   Coefficient 0.09516525
         when "110011100010" => A <= "000111100110110001"; -- Line 13   Column 227   Coefficient 0.11883926
         when "110011100011" => A <= "001001000110101001"; -- Line 13   Column 228   Coefficient 0.14224625
         when "110011100100" => A <= "001010101100000111"; -- Line 13   Column 229   Coefficient 0.16701889
         when "110011100101" => A <= "001100001011101000"; -- Line 13   Column 230   Coefficient 0.19033813
         when "110011100110" => A <= "001101100011111111"; -- Line 13   Column 231   Coefficient 0.21191025
         when "110011100111" => A <= "001110110101010100"; -- Line 13   Column 232   Coefficient 0.23176575
         when "110011101000" => A <= "001111111010100001"; -- Line 13   Column 233   Coefficient 0.24866104
         when "110011101001" => A <= "010000111010100101"; -- Line 13   Column 234   Coefficient 0.26430130
         when "110011101010" => A <= "010010000001100011"; -- Line 13   Column 235   Coefficient 0.28162766
         when "110011101011" => A <= "010010110100110100"; -- Line 13   Column 236   Coefficient 0.29414368
         when "110011101100" => A <= "010011010010100110"; -- Line 13   Column 237   Coefficient 0.30141449
         when "110011101101" => A <= "010011000101100111"; -- Line 13   Column 238   Coefficient 0.29824448
         when "110011101110" => A <= "010001011110001011"; -- Line 13   Column 239   Coefficient 0.27299118
         when "110011101111" => A <= "001111100101110011"; -- Line 13   Column 240   Coefficient 0.24360275
         when "110011110000" => A <= "001101110100101001"; -- Line 13   Column 241   Coefficient 0.21597672
         when "110011110001" => A <= "001011111101111010"; -- Line 13   Column 242   Coefficient 0.18698883
         when "110011110010" => A <= "001010011001111000"; -- Line 13   Column 243   Coefficient 0.16256714
         when "110011110011" => A <= "001000110101000000"; -- Line 13   Column 244   Coefficient 0.13793945
         when "110011110100" => A <= "000111000101010101"; -- Line 13   Column 245   Coefficient 0.11067581
         when "110011110101" => A <= "000101100000010101"; -- Line 13   Column 246   Coefficient 0.08601761
         when "110011110110" => A <= "000100010011001101"; -- Line 13   Column 247   Coefficient 0.06718826
         when "110011110111" => A <= "000011001010010011"; -- Line 13   Column 248   Coefficient 0.04938889
         when "110011111000" => A <= "000010000100001011"; -- Line 13   Column 249   Coefficient 0.03226852
         when "110011111001" => A <= "000000111110100110"; -- Line 13   Column 250   Coefficient 0.01528168
         when "110011111010" => A <= "111111101010001000"; -- Line 13   Column 251   Coefficient -0.00534058
         when "110011111011" => A <= "111110100000101100"; -- Line 13   Column 252   Coefficient -0.02326965
         when "110011111100" => A <= "111101100111001110"; -- Line 13   Column 253   Coefficient -0.03730011
         when "110011111101" => A <= "111101000110110001"; -- Line 13   Column 254   Coefficient -0.04522324
         when "110011111110" => A <= "111101011101101101"; -- Line 13   Column 255   Coefficient -0.03962326
         when "110011111111" => A <= "111101111110110001"; -- Line 13   Column 256   Coefficient -0.03155136
         when "110100000000" => A <= "001101110100101001"; -- Line 14   Column 1   Coefficient 0.21597672
         when "110100000001" => A <= "001011111101111010"; -- Line 14   Column 2   Coefficient 0.18698883
         when "110100000010" => A <= "001010011001111000"; -- Line 14   Column 3   Coefficient 0.16256714
         when "110100000011" => A <= "001000110101000000"; -- Line 14   Column 4   Coefficient 0.13793945
         when "110100000100" => A <= "000111000101010101"; -- Line 14   Column 5   Coefficient 0.11067581
         when "110100000101" => A <= "000101100000010101"; -- Line 14   Column 6   Coefficient 0.08601761
         when "110100000110" => A <= "000100010011001101"; -- Line 14   Column 7   Coefficient 0.06718826
         when "110100000111" => A <= "000011001010010011"; -- Line 14   Column 8   Coefficient 0.04938889
         when "110100001000" => A <= "000010000100001011"; -- Line 14   Column 9   Coefficient 0.03226852
         when "110100001001" => A <= "000000111110100110"; -- Line 14   Column 10   Coefficient 0.01528168
         when "110100001010" => A <= "111111101010001000"; -- Line 14   Column 11   Coefficient -0.00534058
         when "110100001011" => A <= "111110100000101100"; -- Line 14   Column 12   Coefficient -0.02326965
         when "110100001100" => A <= "111101100111001110"; -- Line 14   Column 13   Coefficient -0.03730011
         when "110100001101" => A <= "111101000110110001"; -- Line 14   Column 14   Coefficient -0.04522324
         when "110100001110" => A <= "111101011101101101"; -- Line 14   Column 15   Coefficient -0.03962326
         when "110100001111" => A <= "111101111110110001"; -- Line 14   Column 16   Coefficient -0.03155136
         when "110100010000" => A <= "111110011010010101"; -- Line 14   Column 17   Coefficient -0.02482224
         when "110100010001" => A <= "111110111010000001"; -- Line 14   Column 18   Coefficient -0.01708603
         when "110100010010" => A <= "111111010000101110"; -- Line 14   Column 19   Coefficient -0.01154327
         when "110100010011" => A <= "111111100111100010"; -- Line 14   Column 20   Coefficient -0.00597382
         when "110100010100" => A <= "000000000100100100"; -- Line 14   Column 21   Coefficient 0.00111389
         when "110100010101" => A <= "000000011000110111"; -- Line 14   Column 22   Coefficient 0.00606918
         when "110100010110" => A <= "000000010111101010"; -- Line 14   Column 23   Coefficient 0.00577545
         when "110100010111" => A <= "000000010100111001"; -- Line 14   Column 24   Coefficient 0.00510025
         when "110100011000" => A <= "000000010100110111"; -- Line 14   Column 25   Coefficient 0.00509262
         when "110100011001" => A <= "000000010110010000"; -- Line 14   Column 26   Coefficient 0.00543213
         when "110100011010" => A <= "000000100010100100"; -- Line 14   Column 27   Coefficient 0.00843811
         when "110100011011" => A <= "000000101101010111"; -- Line 14   Column 28   Coefficient 0.01107407
         when "110100011100" => A <= "000000110010101110"; -- Line 14   Column 29   Coefficient 0.01238251
         when "110100011101" => A <= "000000110100010110"; -- Line 14   Column 30   Coefficient 0.01277924
         when "110100011110" => A <= "000000101011110101"; -- Line 14   Column 31   Coefficient 0.01070023
         when "110100011111" => A <= "000000100001110011"; -- Line 14   Column 32   Coefficient 0.00825119
         when "110100100000" => A <= "000000011001110100"; -- Line 14   Column 33   Coefficient 0.00630188
         when "110100100001" => A <= "000000010001001000"; -- Line 14   Column 34   Coefficient 0.00418091
         when "110100100010" => A <= "000000001001011000"; -- Line 14   Column 35   Coefficient 0.00228882
         when "110100100011" => A <= "000000000010010011"; -- Line 14   Column 36   Coefficient 0.00056076
         when "110100100100" => A <= "111111111010111001"; -- Line 14   Column 37   Coefficient -0.00124741
         when "110100100101" => A <= "111111110110011111"; -- Line 14   Column 38   Coefficient -0.00232315
         when "110100100110" => A <= "111111111001000110"; -- Line 14   Column 39   Coefficient -0.00168610
         when "110100100111" => A <= "111111111100011110"; -- Line 14   Column 40   Coefficient -0.00086212
         when "110100101000" => A <= "111111111110110111"; -- Line 14   Column 41   Coefficient -0.00027847
         when "110100101001" => A <= "000000000001001011"; -- Line 14   Column 42   Coefficient 0.00028610
         when "110100101010" => A <= "000000000001001000"; -- Line 14   Column 43   Coefficient 0.00027466
         when "110100101011" => A <= "000000000001000010"; -- Line 14   Column 44   Coefficient 0.00025177
         when "110100101100" => A <= "000000000001111110"; -- Line 14   Column 45   Coefficient 0.00048065
         when "110100101101" => A <= "000000000010010101"; -- Line 14   Column 46   Coefficient 0.00056839
         when "110100101110" => A <= "000000000001100101"; -- Line 14   Column 47   Coefficient 0.00038528
         when "110100101111" => A <= "000000000000110011"; -- Line 14   Column 48   Coefficient 0.00019455
         when "110100110000" => A <= "000000000000000111"; -- Line 14   Column 49   Coefficient 0.00002670
         when "110100110001" => A <= "111111111111100110"; -- Line 14   Column 50   Coefficient -0.00009918
         when "110100110010" => A <= "111111111111110100"; -- Line 14   Column 51   Coefficient -0.00004578
         when "110100110011" => A <= "000000000000000011"; -- Line 14   Column 52   Coefficient 0.00001144
         when "110100110100" => A <= "000000000000000100"; -- Line 14   Column 53   Coefficient 0.00001526
         when "110100110101" => A <= "000000000000000110"; -- Line 14   Column 54   Coefficient 0.00002289
         when "110100110110" => A <= "000000000000000011"; -- Line 14   Column 55   Coefficient 0.00001144
         when "110100110111" => A <= "111111111111111111"; -- Line 14   Column 56   Coefficient -0.00000381
         when "110100111000" => A <= "000000000000000000"; -- Line 14   Column 57   Coefficient 0.00000000
         when "110100111001" => A <= "000000000000000000"; -- Line 14   Column 58   Coefficient 0.00000000
         when "110100111010" => A <= "000000000000000000"; -- Line 14   Column 59   Coefficient 0.00000000
         when "110100111011" => A <= "000000000000000000"; -- Line 14   Column 60   Coefficient 0.00000000
         when "110100111100" => A <= "000000000000000000"; -- Line 14   Column 61   Coefficient 0.00000000
         when "110100111101" => A <= "000000000000000000"; -- Line 14   Column 62   Coefficient 0.00000000
         when "110100111110" => A <= "000000000000000000"; -- Line 14   Column 63   Coefficient 0.00000000
         when "110100111111" => A <= "000000000000000000"; -- Line 14   Column 64   Coefficient 0.00000000
         when "110101000000" => A <= "000000000000000000"; -- Line 14   Column 65   Coefficient 0.00000000
         when "110101000001" => A <= "000000000000000000"; -- Line 14   Column 66   Coefficient 0.00000000
         when "110101000010" => A <= "000000000000000000"; -- Line 14   Column 67   Coefficient 0.00000000
         when "110101000011" => A <= "000000000000000000"; -- Line 14   Column 68   Coefficient 0.00000000
         when "110101000100" => A <= "000000000000000000"; -- Line 14   Column 69   Coefficient 0.00000000
         when "110101000101" => A <= "000000000000000000"; -- Line 14   Column 70   Coefficient 0.00000000
         when "110101000110" => A <= "000000000000000000"; -- Line 14   Column 71   Coefficient 0.00000000
         when "110101000111" => A <= "000000000000000000"; -- Line 14   Column 72   Coefficient 0.00000000
         when "110101001000" => A <= "000000000000000000"; -- Line 14   Column 73   Coefficient 0.00000000
         when "110101001001" => A <= "000000000000000000"; -- Line 14   Column 74   Coefficient 0.00000000
         when "110101001010" => A <= "000000000000000000"; -- Line 14   Column 75   Coefficient 0.00000000
         when "110101001011" => A <= "000000000000000000"; -- Line 14   Column 76   Coefficient 0.00000000
         when "110101001100" => A <= "000000000000000000"; -- Line 14   Column 77   Coefficient 0.00000000
         when "110101001101" => A <= "000000000000000000"; -- Line 14   Column 78   Coefficient 0.00000000
         when "110101001110" => A <= "000000000000000000"; -- Line 14   Column 79   Coefficient 0.00000000
         when "110101001111" => A <= "000000000000000000"; -- Line 14   Column 80   Coefficient 0.00000000
         when "110101010000" => A <= "000000000000000000"; -- Line 14   Column 81   Coefficient 0.00000000
         when "110101010001" => A <= "000000000000000000"; -- Line 14   Column 82   Coefficient 0.00000000
         when "110101010010" => A <= "000000000000000000"; -- Line 14   Column 83   Coefficient 0.00000000
         when "110101010011" => A <= "000000000000000000"; -- Line 14   Column 84   Coefficient 0.00000000
         when "110101010100" => A <= "000000000000000000"; -- Line 14   Column 85   Coefficient 0.00000000
         when "110101010101" => A <= "000000000000000000"; -- Line 14   Column 86   Coefficient 0.00000000
         when "110101010110" => A <= "000000000000000000"; -- Line 14   Column 87   Coefficient 0.00000000
         when "110101010111" => A <= "000000000000000000"; -- Line 14   Column 88   Coefficient 0.00000000
         when "110101011000" => A <= "000000000000000000"; -- Line 14   Column 89   Coefficient 0.00000000
         when "110101011001" => A <= "000000000000000000"; -- Line 14   Column 90   Coefficient 0.00000000
         when "110101011010" => A <= "000000000000000000"; -- Line 14   Column 91   Coefficient 0.00000000
         when "110101011011" => A <= "000000000000000000"; -- Line 14   Column 92   Coefficient 0.00000000
         when "110101011100" => A <= "000000000000000000"; -- Line 14   Column 93   Coefficient 0.00000000
         when "110101011101" => A <= "000000000000000000"; -- Line 14   Column 94   Coefficient 0.00000000
         when "110101011110" => A <= "000000000000000000"; -- Line 14   Column 95   Coefficient 0.00000000
         when "110101011111" => A <= "000000000000000000"; -- Line 14   Column 96   Coefficient 0.00000000
         when "110101100000" => A <= "000000000000000000"; -- Line 14   Column 97   Coefficient 0.00000000
         when "110101100001" => A <= "000000000000000000"; -- Line 14   Column 98   Coefficient 0.00000000
         when "110101100010" => A <= "000000000000000000"; -- Line 14   Column 99   Coefficient 0.00000000
         when "110101100011" => A <= "000000000000000000"; -- Line 14   Column 100   Coefficient 0.00000000
         when "110101100100" => A <= "000000000000000000"; -- Line 14   Column 101   Coefficient 0.00000000
         when "110101100101" => A <= "000000000000000000"; -- Line 14   Column 102   Coefficient 0.00000000
         when "110101100110" => A <= "000000000000000000"; -- Line 14   Column 103   Coefficient 0.00000000
         when "110101100111" => A <= "000000000000000000"; -- Line 14   Column 104   Coefficient 0.00000000
         when "110101101000" => A <= "000000000000000000"; -- Line 14   Column 105   Coefficient 0.00000000
         when "110101101001" => A <= "000000000000000000"; -- Line 14   Column 106   Coefficient 0.00000000
         when "110101101010" => A <= "000000000000000000"; -- Line 14   Column 107   Coefficient 0.00000000
         when "110101101011" => A <= "000000000000000000"; -- Line 14   Column 108   Coefficient 0.00000000
         when "110101101100" => A <= "000000000000000000"; -- Line 14   Column 109   Coefficient 0.00000000
         when "110101101101" => A <= "000000000000000000"; -- Line 14   Column 110   Coefficient 0.00000000
         when "110101101110" => A <= "000000000000000000"; -- Line 14   Column 111   Coefficient 0.00000000
         when "110101101111" => A <= "000000000000000000"; -- Line 14   Column 112   Coefficient 0.00000000
         when "110101110000" => A <= "000000000000000000"; -- Line 14   Column 113   Coefficient 0.00000000
         when "110101110001" => A <= "000000000000000000"; -- Line 14   Column 114   Coefficient 0.00000000
         when "110101110010" => A <= "000000000000000000"; -- Line 14   Column 115   Coefficient 0.00000000
         when "110101110011" => A <= "000000000000000000"; -- Line 14   Column 116   Coefficient 0.00000000
         when "110101110100" => A <= "000000000000000000"; -- Line 14   Column 117   Coefficient 0.00000000
         when "110101110101" => A <= "000000000000000000"; -- Line 14   Column 118   Coefficient 0.00000000
         when "110101110110" => A <= "000000000000000000"; -- Line 14   Column 119   Coefficient 0.00000000
         when "110101110111" => A <= "000000000000000000"; -- Line 14   Column 120   Coefficient 0.00000000
         when "110101111000" => A <= "000000000000000000"; -- Line 14   Column 121   Coefficient 0.00000000
         when "110101111001" => A <= "000000000000000000"; -- Line 14   Column 122   Coefficient 0.00000000
         when "110101111010" => A <= "000000000000000000"; -- Line 14   Column 123   Coefficient 0.00000000
         when "110101111011" => A <= "000000000000000000"; -- Line 14   Column 124   Coefficient 0.00000000
         when "110101111100" => A <= "000000000000000000"; -- Line 14   Column 125   Coefficient 0.00000000
         when "110101111101" => A <= "000000000000000000"; -- Line 14   Column 126   Coefficient 0.00000000
         when "110101111110" => A <= "000000000000000000"; -- Line 14   Column 127   Coefficient 0.00000000
         when "110101111111" => A <= "000000000000000000"; -- Line 14   Column 128   Coefficient 0.00000000
         when "110110000000" => A <= "000000000000000000"; -- Line 14   Column 129   Coefficient 0.00000000
         when "110110000001" => A <= "000000000000000000"; -- Line 14   Column 130   Coefficient 0.00000000
         when "110110000010" => A <= "000000000000000000"; -- Line 14   Column 131   Coefficient 0.00000000
         when "110110000011" => A <= "000000000000000000"; -- Line 14   Column 132   Coefficient 0.00000000
         when "110110000100" => A <= "000000000000000000"; -- Line 14   Column 133   Coefficient 0.00000000
         when "110110000101" => A <= "000000000000000000"; -- Line 14   Column 134   Coefficient 0.00000000
         when "110110000110" => A <= "000000000000000000"; -- Line 14   Column 135   Coefficient 0.00000000
         when "110110000111" => A <= "000000000000000000"; -- Line 14   Column 136   Coefficient 0.00000000
         when "110110001000" => A <= "000000000000000000"; -- Line 14   Column 137   Coefficient 0.00000000
         when "110110001001" => A <= "000000000000000000"; -- Line 14   Column 138   Coefficient 0.00000000
         when "110110001010" => A <= "000000000000000000"; -- Line 14   Column 139   Coefficient 0.00000000
         when "110110001011" => A <= "000000000000000000"; -- Line 14   Column 140   Coefficient 0.00000000
         when "110110001100" => A <= "000000000000000000"; -- Line 14   Column 141   Coefficient 0.00000000
         when "110110001101" => A <= "000000000000000000"; -- Line 14   Column 142   Coefficient 0.00000000
         when "110110001110" => A <= "000000000000000000"; -- Line 14   Column 143   Coefficient 0.00000000
         when "110110001111" => A <= "000000000000000000"; -- Line 14   Column 144   Coefficient 0.00000000
         when "110110010000" => A <= "000000000000000000"; -- Line 14   Column 145   Coefficient 0.00000000
         when "110110010001" => A <= "000000000000000000"; -- Line 14   Column 146   Coefficient 0.00000000
         when "110110010010" => A <= "000000000000000000"; -- Line 14   Column 147   Coefficient 0.00000000
         when "110110010011" => A <= "000000000000000000"; -- Line 14   Column 148   Coefficient 0.00000000
         when "110110010100" => A <= "000000000000000000"; -- Line 14   Column 149   Coefficient 0.00000000
         when "110110010101" => A <= "000000000000000000"; -- Line 14   Column 150   Coefficient 0.00000000
         when "110110010110" => A <= "000000000000000000"; -- Line 14   Column 151   Coefficient 0.00000000
         when "110110010111" => A <= "000000000000000000"; -- Line 14   Column 152   Coefficient 0.00000000
         when "110110011000" => A <= "000000000000000000"; -- Line 14   Column 153   Coefficient 0.00000000
         when "110110011001" => A <= "000000000000000000"; -- Line 14   Column 154   Coefficient 0.00000000
         when "110110011010" => A <= "000000000000000000"; -- Line 14   Column 155   Coefficient 0.00000000
         when "110110011011" => A <= "000000000000000000"; -- Line 14   Column 156   Coefficient 0.00000000
         when "110110011100" => A <= "000000000000000000"; -- Line 14   Column 157   Coefficient 0.00000000
         when "110110011101" => A <= "000000000000000000"; -- Line 14   Column 158   Coefficient 0.00000000
         when "110110011110" => A <= "000000000000000000"; -- Line 14   Column 159   Coefficient 0.00000000
         when "110110011111" => A <= "000000000000000000"; -- Line 14   Column 160   Coefficient 0.00000000
         when "110110100000" => A <= "000000000000000000"; -- Line 14   Column 161   Coefficient 0.00000000
         when "110110100001" => A <= "000000000000000000"; -- Line 14   Column 162   Coefficient 0.00000000
         when "110110100010" => A <= "000000000000000000"; -- Line 14   Column 163   Coefficient 0.00000000
         when "110110100011" => A <= "000000000000000000"; -- Line 14   Column 164   Coefficient 0.00000000
         when "110110100100" => A <= "000000000000000000"; -- Line 14   Column 165   Coefficient 0.00000000
         when "110110100101" => A <= "000000000000000000"; -- Line 14   Column 166   Coefficient 0.00000000
         when "110110100110" => A <= "000000000000000000"; -- Line 14   Column 167   Coefficient 0.00000000
         when "110110100111" => A <= "000000000000000000"; -- Line 14   Column 168   Coefficient 0.00000000
         when "110110101000" => A <= "000000000000000000"; -- Line 14   Column 169   Coefficient 0.00000000
         when "110110101001" => A <= "000000000000000000"; -- Line 14   Column 170   Coefficient 0.00000000
         when "110110101010" => A <= "000000000000000000"; -- Line 14   Column 171   Coefficient 0.00000000
         when "110110101011" => A <= "000000000000000000"; -- Line 14   Column 172   Coefficient 0.00000000
         when "110110101100" => A <= "000000000000000000"; -- Line 14   Column 173   Coefficient 0.00000000
         when "110110101101" => A <= "000000000000000000"; -- Line 14   Column 174   Coefficient 0.00000000
         when "110110101110" => A <= "000000000000000000"; -- Line 14   Column 175   Coefficient 0.00000000
         when "110110101111" => A <= "000000000000000000"; -- Line 14   Column 176   Coefficient 0.00000000
         when "110110110000" => A <= "000000000000000000"; -- Line 14   Column 177   Coefficient 0.00000000
         when "110110110001" => A <= "000000000000000000"; -- Line 14   Column 178   Coefficient 0.00000000
         when "110110110010" => A <= "000000000000000000"; -- Line 14   Column 179   Coefficient 0.00000000
         when "110110110011" => A <= "000000000000000000"; -- Line 14   Column 180   Coefficient 0.00000000
         when "110110110100" => A <= "000000000000000000"; -- Line 14   Column 181   Coefficient 0.00000000
         when "110110110101" => A <= "000000000000000000"; -- Line 14   Column 182   Coefficient 0.00000000
         when "110110110110" => A <= "000000000000000000"; -- Line 14   Column 183   Coefficient 0.00000000
         when "110110110111" => A <= "000000000000000000"; -- Line 14   Column 184   Coefficient 0.00000000
         when "110110111000" => A <= "000000000000000000"; -- Line 14   Column 185   Coefficient 0.00000000
         when "110110111001" => A <= "000000000000000000"; -- Line 14   Column 186   Coefficient 0.00000000
         when "110110111010" => A <= "000000000000000000"; -- Line 14   Column 187   Coefficient 0.00000000
         when "110110111011" => A <= "000000000000000000"; -- Line 14   Column 188   Coefficient 0.00000000
         when "110110111100" => A <= "000000000000000000"; -- Line 14   Column 189   Coefficient 0.00000000
         when "110110111101" => A <= "000000000000000000"; -- Line 14   Column 190   Coefficient 0.00000000
         when "110110111110" => A <= "000000000000000000"; -- Line 14   Column 191   Coefficient 0.00000000
         when "110110111111" => A <= "000000000000000000"; -- Line 14   Column 192   Coefficient 0.00000000
         when "110111000000" => A <= "000000000000000000"; -- Line 14   Column 193   Coefficient 0.00000000
         when "110111000001" => A <= "000000000000000000"; -- Line 14   Column 194   Coefficient 0.00000000
         when "110111000010" => A <= "000000000000000000"; -- Line 14   Column 195   Coefficient 0.00000000
         when "110111000011" => A <= "000000000000000000"; -- Line 14   Column 196   Coefficient 0.00000000
         when "110111000100" => A <= "000000000000000000"; -- Line 14   Column 197   Coefficient 0.00000000
         when "110111000101" => A <= "000000000000000000"; -- Line 14   Column 198   Coefficient 0.00000000
         when "110111000110" => A <= "000000000000000000"; -- Line 14   Column 199   Coefficient 0.00000000
         when "110111000111" => A <= "000000000000000000"; -- Line 14   Column 200   Coefficient 0.00000000
         when "110111001000" => A <= "000000000000000000"; -- Line 14   Column 201   Coefficient 0.00000000
         when "110111001001" => A <= "000000000000000000"; -- Line 14   Column 202   Coefficient 0.00000000
         when "110111001010" => A <= "000000000000000000"; -- Line 14   Column 203   Coefficient 0.00000000
         when "110111001011" => A <= "000000000000000000"; -- Line 14   Column 204   Coefficient 0.00000000
         when "110111001100" => A <= "000000000000000000"; -- Line 14   Column 205   Coefficient 0.00000000
         when "110111001101" => A <= "000000000000000000"; -- Line 14   Column 206   Coefficient 0.00000000
         when "110111001110" => A <= "000000000000000000"; -- Line 14   Column 207   Coefficient 0.00000000
         when "110111001111" => A <= "000000000000000000"; -- Line 14   Column 208   Coefficient 0.00000000
         when "110111010000" => A <= "000000000000001001"; -- Line 14   Column 209   Coefficient 0.00003433
         when "110111010001" => A <= "000000000000000011"; -- Line 14   Column 210   Coefficient 0.00001144
         when "110111010010" => A <= "111111111111001011"; -- Line 14   Column 211   Coefficient -0.00020218
         when "110111010011" => A <= "111111111110100110"; -- Line 14   Column 212   Coefficient -0.00034332
         when "110111010100" => A <= "111111111110010010"; -- Line 14   Column 213   Coefficient -0.00041962
         when "110111010101" => A <= "111111111111010011"; -- Line 14   Column 214   Coefficient -0.00017166
         when "110111010110" => A <= "000000000011111000"; -- Line 14   Column 215   Coefficient 0.00094604
         when "110111010111" => A <= "000000001000010011"; -- Line 14   Column 216   Coefficient 0.00202560
         when "110111011000" => A <= "000000001010110110"; -- Line 14   Column 217   Coefficient 0.00264740
         when "110111011001" => A <= "000000001101001100"; -- Line 14   Column 218   Coefficient 0.00321960
         when "110111011010" => A <= "000000001111111100"; -- Line 14   Column 219   Coefficient 0.00389099
         when "110111011011" => A <= "000000010000011000"; -- Line 14   Column 220   Coefficient 0.00399780
         when "110111011100" => A <= "000000001111000010"; -- Line 14   Column 221   Coefficient 0.00366974
         when "110111011101" => A <= "000000000111011010"; -- Line 14   Column 222   Coefficient 0.00180817
         when "110111011110" => A <= "111111110001010101"; -- Line 14   Column 223   Coefficient -0.00358200
         when "110111011111" => A <= "111111011001111001"; -- Line 14   Column 224   Coefficient -0.00930405
         when "110111100000" => A <= "111111000100111001"; -- Line 14   Column 225   Coefficient -0.01443100
         when "110111100001" => A <= "111110110001100001"; -- Line 14   Column 226   Coefficient -0.01916122
         when "110111100010" => A <= "111110100110010011"; -- Line 14   Column 227   Coefficient -0.02190018
         when "110111100011" => A <= "111110011011111010"; -- Line 14   Column 228   Coefficient -0.02443695
         when "110111100100" => A <= "111110010000110000"; -- Line 14   Column 229   Coefficient -0.02716064
         when "110111100101" => A <= "111110000101010011"; -- Line 14   Column 230   Coefficient -0.02995682
         when "110111100110" => A <= "111101110100001010"; -- Line 14   Column 231   Coefficient -0.03414154
         when "110111100111" => A <= "111101100110110000"; -- Line 14   Column 232   Coefficient -0.03741455
         when "110111101000" => A <= "111101100010101111"; -- Line 14   Column 233   Coefficient -0.03839493
         when "110111101001" => A <= "111101100010001110"; -- Line 14   Column 234   Coefficient -0.03852081
         when "110111101010" => A <= "111101100000101101"; -- Line 14   Column 235   Coefficient -0.03889084
         when "110111101011" => A <= "111101101011101110"; -- Line 14   Column 236   Coefficient -0.03620148
         when "110111101100" => A <= "111110000010011110"; -- Line 14   Column 237   Coefficient -0.03064728
         when "110111101101" => A <= "111110110101100100"; -- Line 14   Column 238   Coefficient -0.01817322
         when "110111101110" => A <= "000000100101011001"; -- Line 14   Column 239   Coefficient 0.00912857
         when "110111101111" => A <= "000010011110111100"; -- Line 14   Column 240   Coefficient 0.03880310
         when "110111110000" => A <= "000100010010000101"; -- Line 14   Column 241   Coefficient 0.06691360
         when "110111110001" => A <= "000110000101110011"; -- Line 14   Column 242   Coefficient 0.09516525
         when "110111110010" => A <= "000111100110110001"; -- Line 14   Column 243   Coefficient 0.11883926
         when "110111110011" => A <= "001001000110101001"; -- Line 14   Column 244   Coefficient 0.14224625
         when "110111110100" => A <= "001010101100000111"; -- Line 14   Column 245   Coefficient 0.16701889
         when "110111110101" => A <= "001100001011101000"; -- Line 14   Column 246   Coefficient 0.19033813
         when "110111110110" => A <= "001101100011111111"; -- Line 14   Column 247   Coefficient 0.21191025
         when "110111110111" => A <= "001110110101010100"; -- Line 14   Column 248   Coefficient 0.23176575
         when "110111111000" => A <= "001111111010100001"; -- Line 14   Column 249   Coefficient 0.24866104
         when "110111111001" => A <= "010000111010100101"; -- Line 14   Column 250   Coefficient 0.26430130
         when "110111111010" => A <= "010010000001100011"; -- Line 14   Column 251   Coefficient 0.28162766
         when "110111111011" => A <= "010010110100110100"; -- Line 14   Column 252   Coefficient 0.29414368
         when "110111111100" => A <= "010011010010100110"; -- Line 14   Column 253   Coefficient 0.30141449
         when "110111111101" => A <= "010011000101100111"; -- Line 14   Column 254   Coefficient 0.29824448
         when "110111111110" => A <= "010001011110001011"; -- Line 14   Column 255   Coefficient 0.27299118
         when "110111111111" => A <= "001111100101110011"; -- Line 14   Column 256   Coefficient 0.24360275
         when "111000000000" => A <= "000100010010000101"; -- Line 15   Column 1   Coefficient 0.06691360
         when "111000000001" => A <= "000110000101110011"; -- Line 15   Column 2   Coefficient 0.09516525
         when "111000000010" => A <= "000111100110110001"; -- Line 15   Column 3   Coefficient 0.11883926
         when "111000000011" => A <= "001001000110101001"; -- Line 15   Column 4   Coefficient 0.14224625
         when "111000000100" => A <= "001010101100000111"; -- Line 15   Column 5   Coefficient 0.16701889
         when "111000000101" => A <= "001100001011101000"; -- Line 15   Column 6   Coefficient 0.19033813
         when "111000000110" => A <= "001101100011111111"; -- Line 15   Column 7   Coefficient 0.21191025
         when "111000000111" => A <= "001110110101010100"; -- Line 15   Column 8   Coefficient 0.23176575
         when "111000001000" => A <= "001111111010100001"; -- Line 15   Column 9   Coefficient 0.24866104
         when "111000001001" => A <= "010000111010100101"; -- Line 15   Column 10   Coefficient 0.26430130
         when "111000001010" => A <= "010010000001100011"; -- Line 15   Column 11   Coefficient 0.28162766
         when "111000001011" => A <= "010010110100110100"; -- Line 15   Column 12   Coefficient 0.29414368
         when "111000001100" => A <= "010011010010100110"; -- Line 15   Column 13   Coefficient 0.30141449
         when "111000001101" => A <= "010011000101100111"; -- Line 15   Column 14   Coefficient 0.29824448
         when "111000001110" => A <= "010001011110001011"; -- Line 15   Column 15   Coefficient 0.27299118
         when "111000001111" => A <= "001111100101110011"; -- Line 15   Column 16   Coefficient 0.24360275
         when "111000010000" => A <= "001101110100101001"; -- Line 15   Column 17   Coefficient 0.21597672
         when "111000010001" => A <= "001011111101111010"; -- Line 15   Column 18   Coefficient 0.18698883
         when "111000010010" => A <= "001010011001111000"; -- Line 15   Column 19   Coefficient 0.16256714
         when "111000010011" => A <= "001000110101000000"; -- Line 15   Column 20   Coefficient 0.13793945
         when "111000010100" => A <= "000111000101010101"; -- Line 15   Column 21   Coefficient 0.11067581
         when "111000010101" => A <= "000101100000010101"; -- Line 15   Column 22   Coefficient 0.08601761
         when "111000010110" => A <= "000100010011001101"; -- Line 15   Column 23   Coefficient 0.06718826
         when "111000010111" => A <= "000011001010010011"; -- Line 15   Column 24   Coefficient 0.04938889
         when "111000011000" => A <= "000010000100001011"; -- Line 15   Column 25   Coefficient 0.03226852
         when "111000011001" => A <= "000000111110100110"; -- Line 15   Column 26   Coefficient 0.01528168
         when "111000011010" => A <= "111111101010001000"; -- Line 15   Column 27   Coefficient -0.00534058
         when "111000011011" => A <= "111110100000101100"; -- Line 15   Column 28   Coefficient -0.02326965
         when "111000011100" => A <= "111101100111001110"; -- Line 15   Column 29   Coefficient -0.03730011
         when "111000011101" => A <= "111101000110110001"; -- Line 15   Column 30   Coefficient -0.04522324
         when "111000011110" => A <= "111101011101101101"; -- Line 15   Column 31   Coefficient -0.03962326
         when "111000011111" => A <= "111101111110110001"; -- Line 15   Column 32   Coefficient -0.03155136
         when "111000100000" => A <= "111110011010010101"; -- Line 15   Column 33   Coefficient -0.02482224
         when "111000100001" => A <= "111110111010000001"; -- Line 15   Column 34   Coefficient -0.01708603
         when "111000100010" => A <= "111111010000101110"; -- Line 15   Column 35   Coefficient -0.01154327
         when "111000100011" => A <= "111111100111100010"; -- Line 15   Column 36   Coefficient -0.00597382
         when "111000100100" => A <= "000000000100100100"; -- Line 15   Column 37   Coefficient 0.00111389
         when "111000100101" => A <= "000000011000110111"; -- Line 15   Column 38   Coefficient 0.00606918
         when "111000100110" => A <= "000000010111101010"; -- Line 15   Column 39   Coefficient 0.00577545
         when "111000100111" => A <= "000000010100111001"; -- Line 15   Column 40   Coefficient 0.00510025
         when "111000101000" => A <= "000000010100110111"; -- Line 15   Column 41   Coefficient 0.00509262
         when "111000101001" => A <= "000000010110010000"; -- Line 15   Column 42   Coefficient 0.00543213
         when "111000101010" => A <= "000000100010100100"; -- Line 15   Column 43   Coefficient 0.00843811
         when "111000101011" => A <= "000000101101010111"; -- Line 15   Column 44   Coefficient 0.01107407
         when "111000101100" => A <= "000000110010101110"; -- Line 15   Column 45   Coefficient 0.01238251
         when "111000101101" => A <= "000000110100010110"; -- Line 15   Column 46   Coefficient 0.01277924
         when "111000101110" => A <= "000000101011110101"; -- Line 15   Column 47   Coefficient 0.01070023
         when "111000101111" => A <= "000000100001110011"; -- Line 15   Column 48   Coefficient 0.00825119
         when "111000110000" => A <= "000000011001110100"; -- Line 15   Column 49   Coefficient 0.00630188
         when "111000110001" => A <= "000000010001001000"; -- Line 15   Column 50   Coefficient 0.00418091
         when "111000110010" => A <= "000000001001011000"; -- Line 15   Column 51   Coefficient 0.00228882
         when "111000110011" => A <= "000000000010010011"; -- Line 15   Column 52   Coefficient 0.00056076
         when "111000110100" => A <= "111111111010111001"; -- Line 15   Column 53   Coefficient -0.00124741
         when "111000110101" => A <= "111111110110011111"; -- Line 15   Column 54   Coefficient -0.00232315
         when "111000110110" => A <= "111111111001000110"; -- Line 15   Column 55   Coefficient -0.00168610
         when "111000110111" => A <= "111111111100011110"; -- Line 15   Column 56   Coefficient -0.00086212
         when "111000111000" => A <= "111111111110110111"; -- Line 15   Column 57   Coefficient -0.00027847
         when "111000111001" => A <= "000000000001001011"; -- Line 15   Column 58   Coefficient 0.00028610
         when "111000111010" => A <= "000000000001001000"; -- Line 15   Column 59   Coefficient 0.00027466
         when "111000111011" => A <= "000000000001000010"; -- Line 15   Column 60   Coefficient 0.00025177
         when "111000111100" => A <= "000000000001111110"; -- Line 15   Column 61   Coefficient 0.00048065
         when "111000111101" => A <= "000000000010010101"; -- Line 15   Column 62   Coefficient 0.00056839
         when "111000111110" => A <= "000000000001100101"; -- Line 15   Column 63   Coefficient 0.00038528
         when "111000111111" => A <= "000000000000110011"; -- Line 15   Column 64   Coefficient 0.00019455
         when "111001000000" => A <= "000000000000000111"; -- Line 15   Column 65   Coefficient 0.00002670
         when "111001000001" => A <= "111111111111100110"; -- Line 15   Column 66   Coefficient -0.00009918
         when "111001000010" => A <= "111111111111110100"; -- Line 15   Column 67   Coefficient -0.00004578
         when "111001000011" => A <= "000000000000000011"; -- Line 15   Column 68   Coefficient 0.00001144
         when "111001000100" => A <= "000000000000000100"; -- Line 15   Column 69   Coefficient 0.00001526
         when "111001000101" => A <= "000000000000000110"; -- Line 15   Column 70   Coefficient 0.00002289
         when "111001000110" => A <= "000000000000000011"; -- Line 15   Column 71   Coefficient 0.00001144
         when "111001000111" => A <= "111111111111111111"; -- Line 15   Column 72   Coefficient -0.00000381
         when "111001001000" => A <= "000000000000000000"; -- Line 15   Column 73   Coefficient 0.00000000
         when "111001001001" => A <= "000000000000000000"; -- Line 15   Column 74   Coefficient 0.00000000
         when "111001001010" => A <= "000000000000000000"; -- Line 15   Column 75   Coefficient 0.00000000
         when "111001001011" => A <= "000000000000000000"; -- Line 15   Column 76   Coefficient 0.00000000
         when "111001001100" => A <= "000000000000000000"; -- Line 15   Column 77   Coefficient 0.00000000
         when "111001001101" => A <= "000000000000000000"; -- Line 15   Column 78   Coefficient 0.00000000
         when "111001001110" => A <= "000000000000000000"; -- Line 15   Column 79   Coefficient 0.00000000
         when "111001001111" => A <= "000000000000000000"; -- Line 15   Column 80   Coefficient 0.00000000
         when "111001010000" => A <= "000000000000000000"; -- Line 15   Column 81   Coefficient 0.00000000
         when "111001010001" => A <= "000000000000000000"; -- Line 15   Column 82   Coefficient 0.00000000
         when "111001010010" => A <= "000000000000000000"; -- Line 15   Column 83   Coefficient 0.00000000
         when "111001010011" => A <= "000000000000000000"; -- Line 15   Column 84   Coefficient 0.00000000
         when "111001010100" => A <= "000000000000000000"; -- Line 15   Column 85   Coefficient 0.00000000
         when "111001010101" => A <= "000000000000000000"; -- Line 15   Column 86   Coefficient 0.00000000
         when "111001010110" => A <= "000000000000000000"; -- Line 15   Column 87   Coefficient 0.00000000
         when "111001010111" => A <= "000000000000000000"; -- Line 15   Column 88   Coefficient 0.00000000
         when "111001011000" => A <= "000000000000000000"; -- Line 15   Column 89   Coefficient 0.00000000
         when "111001011001" => A <= "000000000000000000"; -- Line 15   Column 90   Coefficient 0.00000000
         when "111001011010" => A <= "000000000000000000"; -- Line 15   Column 91   Coefficient 0.00000000
         when "111001011011" => A <= "000000000000000000"; -- Line 15   Column 92   Coefficient 0.00000000
         when "111001011100" => A <= "000000000000000000"; -- Line 15   Column 93   Coefficient 0.00000000
         when "111001011101" => A <= "000000000000000000"; -- Line 15   Column 94   Coefficient 0.00000000
         when "111001011110" => A <= "000000000000000000"; -- Line 15   Column 95   Coefficient 0.00000000
         when "111001011111" => A <= "000000000000000000"; -- Line 15   Column 96   Coefficient 0.00000000
         when "111001100000" => A <= "000000000000000000"; -- Line 15   Column 97   Coefficient 0.00000000
         when "111001100001" => A <= "000000000000000000"; -- Line 15   Column 98   Coefficient 0.00000000
         when "111001100010" => A <= "000000000000000000"; -- Line 15   Column 99   Coefficient 0.00000000
         when "111001100011" => A <= "000000000000000000"; -- Line 15   Column 100   Coefficient 0.00000000
         when "111001100100" => A <= "000000000000000000"; -- Line 15   Column 101   Coefficient 0.00000000
         when "111001100101" => A <= "000000000000000000"; -- Line 15   Column 102   Coefficient 0.00000000
         when "111001100110" => A <= "000000000000000000"; -- Line 15   Column 103   Coefficient 0.00000000
         when "111001100111" => A <= "000000000000000000"; -- Line 15   Column 104   Coefficient 0.00000000
         when "111001101000" => A <= "000000000000000000"; -- Line 15   Column 105   Coefficient 0.00000000
         when "111001101001" => A <= "000000000000000000"; -- Line 15   Column 106   Coefficient 0.00000000
         when "111001101010" => A <= "000000000000000000"; -- Line 15   Column 107   Coefficient 0.00000000
         when "111001101011" => A <= "000000000000000000"; -- Line 15   Column 108   Coefficient 0.00000000
         when "111001101100" => A <= "000000000000000000"; -- Line 15   Column 109   Coefficient 0.00000000
         when "111001101101" => A <= "000000000000000000"; -- Line 15   Column 110   Coefficient 0.00000000
         when "111001101110" => A <= "000000000000000000"; -- Line 15   Column 111   Coefficient 0.00000000
         when "111001101111" => A <= "000000000000000000"; -- Line 15   Column 112   Coefficient 0.00000000
         when "111001110000" => A <= "000000000000000000"; -- Line 15   Column 113   Coefficient 0.00000000
         when "111001110001" => A <= "000000000000000000"; -- Line 15   Column 114   Coefficient 0.00000000
         when "111001110010" => A <= "000000000000000000"; -- Line 15   Column 115   Coefficient 0.00000000
         when "111001110011" => A <= "000000000000000000"; -- Line 15   Column 116   Coefficient 0.00000000
         when "111001110100" => A <= "000000000000000000"; -- Line 15   Column 117   Coefficient 0.00000000
         when "111001110101" => A <= "000000000000000000"; -- Line 15   Column 118   Coefficient 0.00000000
         when "111001110110" => A <= "000000000000000000"; -- Line 15   Column 119   Coefficient 0.00000000
         when "111001110111" => A <= "000000000000000000"; -- Line 15   Column 120   Coefficient 0.00000000
         when "111001111000" => A <= "000000000000000000"; -- Line 15   Column 121   Coefficient 0.00000000
         when "111001111001" => A <= "000000000000000000"; -- Line 15   Column 122   Coefficient 0.00000000
         when "111001111010" => A <= "000000000000000000"; -- Line 15   Column 123   Coefficient 0.00000000
         when "111001111011" => A <= "000000000000000000"; -- Line 15   Column 124   Coefficient 0.00000000
         when "111001111100" => A <= "000000000000000000"; -- Line 15   Column 125   Coefficient 0.00000000
         when "111001111101" => A <= "000000000000000000"; -- Line 15   Column 126   Coefficient 0.00000000
         when "111001111110" => A <= "000000000000000000"; -- Line 15   Column 127   Coefficient 0.00000000
         when "111001111111" => A <= "000000000000000000"; -- Line 15   Column 128   Coefficient 0.00000000
         when "111010000000" => A <= "000000000000000000"; -- Line 15   Column 129   Coefficient 0.00000000
         when "111010000001" => A <= "000000000000000000"; -- Line 15   Column 130   Coefficient 0.00000000
         when "111010000010" => A <= "000000000000000000"; -- Line 15   Column 131   Coefficient 0.00000000
         when "111010000011" => A <= "000000000000000000"; -- Line 15   Column 132   Coefficient 0.00000000
         when "111010000100" => A <= "000000000000000000"; -- Line 15   Column 133   Coefficient 0.00000000
         when "111010000101" => A <= "000000000000000000"; -- Line 15   Column 134   Coefficient 0.00000000
         when "111010000110" => A <= "000000000000000000"; -- Line 15   Column 135   Coefficient 0.00000000
         when "111010000111" => A <= "000000000000000000"; -- Line 15   Column 136   Coefficient 0.00000000
         when "111010001000" => A <= "000000000000000000"; -- Line 15   Column 137   Coefficient 0.00000000
         when "111010001001" => A <= "000000000000000000"; -- Line 15   Column 138   Coefficient 0.00000000
         when "111010001010" => A <= "000000000000000000"; -- Line 15   Column 139   Coefficient 0.00000000
         when "111010001011" => A <= "000000000000000000"; -- Line 15   Column 140   Coefficient 0.00000000
         when "111010001100" => A <= "000000000000000000"; -- Line 15   Column 141   Coefficient 0.00000000
         when "111010001101" => A <= "000000000000000000"; -- Line 15   Column 142   Coefficient 0.00000000
         when "111010001110" => A <= "000000000000000000"; -- Line 15   Column 143   Coefficient 0.00000000
         when "111010001111" => A <= "000000000000000000"; -- Line 15   Column 144   Coefficient 0.00000000
         when "111010010000" => A <= "000000000000000000"; -- Line 15   Column 145   Coefficient 0.00000000
         when "111010010001" => A <= "000000000000000000"; -- Line 15   Column 146   Coefficient 0.00000000
         when "111010010010" => A <= "000000000000000000"; -- Line 15   Column 147   Coefficient 0.00000000
         when "111010010011" => A <= "000000000000000000"; -- Line 15   Column 148   Coefficient 0.00000000
         when "111010010100" => A <= "000000000000000000"; -- Line 15   Column 149   Coefficient 0.00000000
         when "111010010101" => A <= "000000000000000000"; -- Line 15   Column 150   Coefficient 0.00000000
         when "111010010110" => A <= "000000000000000000"; -- Line 15   Column 151   Coefficient 0.00000000
         when "111010010111" => A <= "000000000000000000"; -- Line 15   Column 152   Coefficient 0.00000000
         when "111010011000" => A <= "000000000000000000"; -- Line 15   Column 153   Coefficient 0.00000000
         when "111010011001" => A <= "000000000000000000"; -- Line 15   Column 154   Coefficient 0.00000000
         when "111010011010" => A <= "000000000000000000"; -- Line 15   Column 155   Coefficient 0.00000000
         when "111010011011" => A <= "000000000000000000"; -- Line 15   Column 156   Coefficient 0.00000000
         when "111010011100" => A <= "000000000000000000"; -- Line 15   Column 157   Coefficient 0.00000000
         when "111010011101" => A <= "000000000000000000"; -- Line 15   Column 158   Coefficient 0.00000000
         when "111010011110" => A <= "000000000000000000"; -- Line 15   Column 159   Coefficient 0.00000000
         when "111010011111" => A <= "000000000000000000"; -- Line 15   Column 160   Coefficient 0.00000000
         when "111010100000" => A <= "000000000000000000"; -- Line 15   Column 161   Coefficient 0.00000000
         when "111010100001" => A <= "000000000000000000"; -- Line 15   Column 162   Coefficient 0.00000000
         when "111010100010" => A <= "000000000000000000"; -- Line 15   Column 163   Coefficient 0.00000000
         when "111010100011" => A <= "000000000000000000"; -- Line 15   Column 164   Coefficient 0.00000000
         when "111010100100" => A <= "000000000000000000"; -- Line 15   Column 165   Coefficient 0.00000000
         when "111010100101" => A <= "000000000000000000"; -- Line 15   Column 166   Coefficient 0.00000000
         when "111010100110" => A <= "000000000000000000"; -- Line 15   Column 167   Coefficient 0.00000000
         when "111010100111" => A <= "000000000000000000"; -- Line 15   Column 168   Coefficient 0.00000000
         when "111010101000" => A <= "000000000000000000"; -- Line 15   Column 169   Coefficient 0.00000000
         when "111010101001" => A <= "000000000000000000"; -- Line 15   Column 170   Coefficient 0.00000000
         when "111010101010" => A <= "000000000000000000"; -- Line 15   Column 171   Coefficient 0.00000000
         when "111010101011" => A <= "000000000000000000"; -- Line 15   Column 172   Coefficient 0.00000000
         when "111010101100" => A <= "000000000000000000"; -- Line 15   Column 173   Coefficient 0.00000000
         when "111010101101" => A <= "000000000000000000"; -- Line 15   Column 174   Coefficient 0.00000000
         when "111010101110" => A <= "000000000000000000"; -- Line 15   Column 175   Coefficient 0.00000000
         when "111010101111" => A <= "000000000000000000"; -- Line 15   Column 176   Coefficient 0.00000000
         when "111010110000" => A <= "000000000000000000"; -- Line 15   Column 177   Coefficient 0.00000000
         when "111010110001" => A <= "000000000000000000"; -- Line 15   Column 178   Coefficient 0.00000000
         when "111010110010" => A <= "000000000000000000"; -- Line 15   Column 179   Coefficient 0.00000000
         when "111010110011" => A <= "000000000000000000"; -- Line 15   Column 180   Coefficient 0.00000000
         when "111010110100" => A <= "000000000000000000"; -- Line 15   Column 181   Coefficient 0.00000000
         when "111010110101" => A <= "000000000000000000"; -- Line 15   Column 182   Coefficient 0.00000000
         when "111010110110" => A <= "000000000000000000"; -- Line 15   Column 183   Coefficient 0.00000000
         when "111010110111" => A <= "000000000000000000"; -- Line 15   Column 184   Coefficient 0.00000000
         when "111010111000" => A <= "000000000000000000"; -- Line 15   Column 185   Coefficient 0.00000000
         when "111010111001" => A <= "000000000000000000"; -- Line 15   Column 186   Coefficient 0.00000000
         when "111010111010" => A <= "000000000000000000"; -- Line 15   Column 187   Coefficient 0.00000000
         when "111010111011" => A <= "000000000000000000"; -- Line 15   Column 188   Coefficient 0.00000000
         when "111010111100" => A <= "000000000000000000"; -- Line 15   Column 189   Coefficient 0.00000000
         when "111010111101" => A <= "000000000000000000"; -- Line 15   Column 190   Coefficient 0.00000000
         when "111010111110" => A <= "000000000000000000"; -- Line 15   Column 191   Coefficient 0.00000000
         when "111010111111" => A <= "000000000000000000"; -- Line 15   Column 192   Coefficient 0.00000000
         when "111011000000" => A <= "000000000000000000"; -- Line 15   Column 193   Coefficient 0.00000000
         when "111011000001" => A <= "000000000000000000"; -- Line 15   Column 194   Coefficient 0.00000000
         when "111011000010" => A <= "000000000000000000"; -- Line 15   Column 195   Coefficient 0.00000000
         when "111011000011" => A <= "000000000000000000"; -- Line 15   Column 196   Coefficient 0.00000000
         when "111011000100" => A <= "000000000000000000"; -- Line 15   Column 197   Coefficient 0.00000000
         when "111011000101" => A <= "000000000000000000"; -- Line 15   Column 198   Coefficient 0.00000000
         when "111011000110" => A <= "000000000000000000"; -- Line 15   Column 199   Coefficient 0.00000000
         when "111011000111" => A <= "000000000000000000"; -- Line 15   Column 200   Coefficient 0.00000000
         when "111011001000" => A <= "000000000000000000"; -- Line 15   Column 201   Coefficient 0.00000000
         when "111011001001" => A <= "000000000000000000"; -- Line 15   Column 202   Coefficient 0.00000000
         when "111011001010" => A <= "000000000000000000"; -- Line 15   Column 203   Coefficient 0.00000000
         when "111011001011" => A <= "000000000000000000"; -- Line 15   Column 204   Coefficient 0.00000000
         when "111011001100" => A <= "000000000000000000"; -- Line 15   Column 205   Coefficient 0.00000000
         when "111011001101" => A <= "000000000000000000"; -- Line 15   Column 206   Coefficient 0.00000000
         when "111011001110" => A <= "000000000000000000"; -- Line 15   Column 207   Coefficient 0.00000000
         when "111011001111" => A <= "000000000000000000"; -- Line 15   Column 208   Coefficient 0.00000000
         when "111011010000" => A <= "000000000000000000"; -- Line 15   Column 209   Coefficient 0.00000000
         when "111011010001" => A <= "000000000000000000"; -- Line 15   Column 210   Coefficient 0.00000000
         when "111011010010" => A <= "000000000000000000"; -- Line 15   Column 211   Coefficient 0.00000000
         when "111011010011" => A <= "000000000000000000"; -- Line 15   Column 212   Coefficient 0.00000000
         when "111011010100" => A <= "000000000000000000"; -- Line 15   Column 213   Coefficient 0.00000000
         when "111011010101" => A <= "000000000000000000"; -- Line 15   Column 214   Coefficient 0.00000000
         when "111011010110" => A <= "000000000000000000"; -- Line 15   Column 215   Coefficient 0.00000000
         when "111011010111" => A <= "000000000000000000"; -- Line 15   Column 216   Coefficient 0.00000000
         when "111011011000" => A <= "000000000000000000"; -- Line 15   Column 217   Coefficient 0.00000000
         when "111011011001" => A <= "000000000000000000"; -- Line 15   Column 218   Coefficient 0.00000000
         when "111011011010" => A <= "000000000000000000"; -- Line 15   Column 219   Coefficient 0.00000000
         when "111011011011" => A <= "000000000000000000"; -- Line 15   Column 220   Coefficient 0.00000000
         when "111011011100" => A <= "000000000000000000"; -- Line 15   Column 221   Coefficient 0.00000000
         when "111011011101" => A <= "000000000000000000"; -- Line 15   Column 222   Coefficient 0.00000000
         when "111011011110" => A <= "000000000000000000"; -- Line 15   Column 223   Coefficient 0.00000000
         when "111011011111" => A <= "000000000000000000"; -- Line 15   Column 224   Coefficient 0.00000000
         when "111011100000" => A <= "000000000000001001"; -- Line 15   Column 225   Coefficient 0.00003433
         when "111011100001" => A <= "000000000000000011"; -- Line 15   Column 226   Coefficient 0.00001144
         when "111011100010" => A <= "111111111111001011"; -- Line 15   Column 227   Coefficient -0.00020218
         when "111011100011" => A <= "111111111110100110"; -- Line 15   Column 228   Coefficient -0.00034332
         when "111011100100" => A <= "111111111110010010"; -- Line 15   Column 229   Coefficient -0.00041962
         when "111011100101" => A <= "111111111111010011"; -- Line 15   Column 230   Coefficient -0.00017166
         when "111011100110" => A <= "000000000011111000"; -- Line 15   Column 231   Coefficient 0.00094604
         when "111011100111" => A <= "000000001000010011"; -- Line 15   Column 232   Coefficient 0.00202560
         when "111011101000" => A <= "000000001010110110"; -- Line 15   Column 233   Coefficient 0.00264740
         when "111011101001" => A <= "000000001101001100"; -- Line 15   Column 234   Coefficient 0.00321960
         when "111011101010" => A <= "000000001111111100"; -- Line 15   Column 235   Coefficient 0.00389099
         when "111011101011" => A <= "000000010000011000"; -- Line 15   Column 236   Coefficient 0.00399780
         when "111011101100" => A <= "000000001111000010"; -- Line 15   Column 237   Coefficient 0.00366974
         when "111011101101" => A <= "000000000111011010"; -- Line 15   Column 238   Coefficient 0.00180817
         when "111011101110" => A <= "111111110001010101"; -- Line 15   Column 239   Coefficient -0.00358200
         when "111011101111" => A <= "111111011001111001"; -- Line 15   Column 240   Coefficient -0.00930405
         when "111011110000" => A <= "111111000100111001"; -- Line 15   Column 241   Coefficient -0.01443100
         when "111011110001" => A <= "111110110001100001"; -- Line 15   Column 242   Coefficient -0.01916122
         when "111011110010" => A <= "111110100110010011"; -- Line 15   Column 243   Coefficient -0.02190018
         when "111011110011" => A <= "111110011011111010"; -- Line 15   Column 244   Coefficient -0.02443695
         when "111011110100" => A <= "111110010000110000"; -- Line 15   Column 245   Coefficient -0.02716064
         when "111011110101" => A <= "111110000101010011"; -- Line 15   Column 246   Coefficient -0.02995682
         when "111011110110" => A <= "111101110100001010"; -- Line 15   Column 247   Coefficient -0.03414154
         when "111011110111" => A <= "111101100110110000"; -- Line 15   Column 248   Coefficient -0.03741455
         when "111011111000" => A <= "111101100010101111"; -- Line 15   Column 249   Coefficient -0.03839493
         when "111011111001" => A <= "111101100010001110"; -- Line 15   Column 250   Coefficient -0.03852081
         when "111011111010" => A <= "111101100000101101"; -- Line 15   Column 251   Coefficient -0.03889084
         when "111011111011" => A <= "111101101011101110"; -- Line 15   Column 252   Coefficient -0.03620148
         when "111011111100" => A <= "111110000010011110"; -- Line 15   Column 253   Coefficient -0.03064728
         when "111011111101" => A <= "111110110101100100"; -- Line 15   Column 254   Coefficient -0.01817322
         when "111011111110" => A <= "000000100101011001"; -- Line 15   Column 255   Coefficient 0.00912857
         when "111011111111" => A <= "000010011110111100"; -- Line 15   Column 256   Coefficient 0.03880310
         when "111100000000" => A <= "111111000100111001"; -- Line 16   Column 1   Coefficient -0.01443100
         when "111100000001" => A <= "111110110001100001"; -- Line 16   Column 2   Coefficient -0.01916122
         when "111100000010" => A <= "111110100110010011"; -- Line 16   Column 3   Coefficient -0.02190018
         when "111100000011" => A <= "111110011011111010"; -- Line 16   Column 4   Coefficient -0.02443695
         when "111100000100" => A <= "111110010000110000"; -- Line 16   Column 5   Coefficient -0.02716064
         when "111100000101" => A <= "111110000101010011"; -- Line 16   Column 6   Coefficient -0.02995682
         when "111100000110" => A <= "111101110100001010"; -- Line 16   Column 7   Coefficient -0.03414154
         when "111100000111" => A <= "111101100110110000"; -- Line 16   Column 8   Coefficient -0.03741455
         when "111100001000" => A <= "111101100010101111"; -- Line 16   Column 9   Coefficient -0.03839493
         when "111100001001" => A <= "111101100010001110"; -- Line 16   Column 10   Coefficient -0.03852081
         when "111100001010" => A <= "111101100000101101"; -- Line 16   Column 11   Coefficient -0.03889084
         when "111100001011" => A <= "111101101011101110"; -- Line 16   Column 12   Coefficient -0.03620148
         when "111100001100" => A <= "111110000010011110"; -- Line 16   Column 13   Coefficient -0.03064728
         when "111100001101" => A <= "111110110101100100"; -- Line 16   Column 14   Coefficient -0.01817322
         when "111100001110" => A <= "000000100101011001"; -- Line 16   Column 15   Coefficient 0.00912857
         when "111100001111" => A <= "000010011110111100"; -- Line 16   Column 16   Coefficient 0.03880310
         when "111100010000" => A <= "000100010010000101"; -- Line 16   Column 17   Coefficient 0.06691360
         when "111100010001" => A <= "000110000101110011"; -- Line 16   Column 18   Coefficient 0.09516525
         when "111100010010" => A <= "000111100110110001"; -- Line 16   Column 19   Coefficient 0.11883926
         when "111100010011" => A <= "001001000110101001"; -- Line 16   Column 20   Coefficient 0.14224625
         when "111100010100" => A <= "001010101100000111"; -- Line 16   Column 21   Coefficient 0.16701889
         when "111100010101" => A <= "001100001011101000"; -- Line 16   Column 22   Coefficient 0.19033813
         when "111100010110" => A <= "001101100011111111"; -- Line 16   Column 23   Coefficient 0.21191025
         when "111100010111" => A <= "001110110101010100"; -- Line 16   Column 24   Coefficient 0.23176575
         when "111100011000" => A <= "001111111010100001"; -- Line 16   Column 25   Coefficient 0.24866104
         when "111100011001" => A <= "010000111010100101"; -- Line 16   Column 26   Coefficient 0.26430130
         when "111100011010" => A <= "010010000001100011"; -- Line 16   Column 27   Coefficient 0.28162766
         when "111100011011" => A <= "010010110100110100"; -- Line 16   Column 28   Coefficient 0.29414368
         when "111100011100" => A <= "010011010010100110"; -- Line 16   Column 29   Coefficient 0.30141449
         when "111100011101" => A <= "010011000101100111"; -- Line 16   Column 30   Coefficient 0.29824448
         when "111100011110" => A <= "010001011110001011"; -- Line 16   Column 31   Coefficient 0.27299118
         when "111100011111" => A <= "001111100101110011"; -- Line 16   Column 32   Coefficient 0.24360275
         when "111100100000" => A <= "001101110100101001"; -- Line 16   Column 33   Coefficient 0.21597672
         when "111100100001" => A <= "001011111101111010"; -- Line 16   Column 34   Coefficient 0.18698883
         when "111100100010" => A <= "001010011001111000"; -- Line 16   Column 35   Coefficient 0.16256714
         when "111100100011" => A <= "001000110101000000"; -- Line 16   Column 36   Coefficient 0.13793945
         when "111100100100" => A <= "000111000101010101"; -- Line 16   Column 37   Coefficient 0.11067581
         when "111100100101" => A <= "000101100000010101"; -- Line 16   Column 38   Coefficient 0.08601761
         when "111100100110" => A <= "000100010011001101"; -- Line 16   Column 39   Coefficient 0.06718826
         when "111100100111" => A <= "000011001010010011"; -- Line 16   Column 40   Coefficient 0.04938889
         when "111100101000" => A <= "000010000100001011"; -- Line 16   Column 41   Coefficient 0.03226852
         when "111100101001" => A <= "000000111110100110"; -- Line 16   Column 42   Coefficient 0.01528168
         when "111100101010" => A <= "111111101010001000"; -- Line 16   Column 43   Coefficient -0.00534058
         when "111100101011" => A <= "111110100000101100"; -- Line 16   Column 44   Coefficient -0.02326965
         when "111100101100" => A <= "111101100111001110"; -- Line 16   Column 45   Coefficient -0.03730011
         when "111100101101" => A <= "111101000110110001"; -- Line 16   Column 46   Coefficient -0.04522324
         when "111100101110" => A <= "111101011101101101"; -- Line 16   Column 47   Coefficient -0.03962326
         when "111100101111" => A <= "111101111110110001"; -- Line 16   Column 48   Coefficient -0.03155136
         when "111100110000" => A <= "111110011010010101"; -- Line 16   Column 49   Coefficient -0.02482224
         when "111100110001" => A <= "111110111010000001"; -- Line 16   Column 50   Coefficient -0.01708603
         when "111100110010" => A <= "111111010000101110"; -- Line 16   Column 51   Coefficient -0.01154327
         when "111100110011" => A <= "111111100111100010"; -- Line 16   Column 52   Coefficient -0.00597382
         when "111100110100" => A <= "000000000100100100"; -- Line 16   Column 53   Coefficient 0.00111389
         when "111100110101" => A <= "000000011000110111"; -- Line 16   Column 54   Coefficient 0.00606918
         when "111100110110" => A <= "000000010111101010"; -- Line 16   Column 55   Coefficient 0.00577545
         when "111100110111" => A <= "000000010100111001"; -- Line 16   Column 56   Coefficient 0.00510025
         when "111100111000" => A <= "000000010100110111"; -- Line 16   Column 57   Coefficient 0.00509262
         when "111100111001" => A <= "000000010110010000"; -- Line 16   Column 58   Coefficient 0.00543213
         when "111100111010" => A <= "000000100010100100"; -- Line 16   Column 59   Coefficient 0.00843811
         when "111100111011" => A <= "000000101101010111"; -- Line 16   Column 60   Coefficient 0.01107407
         when "111100111100" => A <= "000000110010101110"; -- Line 16   Column 61   Coefficient 0.01238251
         when "111100111101" => A <= "000000110100010110"; -- Line 16   Column 62   Coefficient 0.01277924
         when "111100111110" => A <= "000000101011110101"; -- Line 16   Column 63   Coefficient 0.01070023
         when "111100111111" => A <= "000000100001110011"; -- Line 16   Column 64   Coefficient 0.00825119
         when "111101000000" => A <= "000000011001110100"; -- Line 16   Column 65   Coefficient 0.00630188
         when "111101000001" => A <= "000000010001001000"; -- Line 16   Column 66   Coefficient 0.00418091
         when "111101000010" => A <= "000000001001011000"; -- Line 16   Column 67   Coefficient 0.00228882
         when "111101000011" => A <= "000000000010010011"; -- Line 16   Column 68   Coefficient 0.00056076
         when "111101000100" => A <= "111111111010111001"; -- Line 16   Column 69   Coefficient -0.00124741
         when "111101000101" => A <= "111111110110011111"; -- Line 16   Column 70   Coefficient -0.00232315
         when "111101000110" => A <= "111111111001000110"; -- Line 16   Column 71   Coefficient -0.00168610
         when "111101000111" => A <= "111111111100011110"; -- Line 16   Column 72   Coefficient -0.00086212
         when "111101001000" => A <= "111111111110110111"; -- Line 16   Column 73   Coefficient -0.00027847
         when "111101001001" => A <= "000000000001001011"; -- Line 16   Column 74   Coefficient 0.00028610
         when "111101001010" => A <= "000000000001001000"; -- Line 16   Column 75   Coefficient 0.00027466
         when "111101001011" => A <= "000000000001000010"; -- Line 16   Column 76   Coefficient 0.00025177
         when "111101001100" => A <= "000000000001111110"; -- Line 16   Column 77   Coefficient 0.00048065
         when "111101001101" => A <= "000000000010010101"; -- Line 16   Column 78   Coefficient 0.00056839
         when "111101001110" => A <= "000000000001100101"; -- Line 16   Column 79   Coefficient 0.00038528
         when "111101001111" => A <= "000000000000110011"; -- Line 16   Column 80   Coefficient 0.00019455
         when "111101010000" => A <= "000000000000000111"; -- Line 16   Column 81   Coefficient 0.00002670
         when "111101010001" => A <= "111111111111100110"; -- Line 16   Column 82   Coefficient -0.00009918
         when "111101010010" => A <= "111111111111110100"; -- Line 16   Column 83   Coefficient -0.00004578
         when "111101010011" => A <= "000000000000000011"; -- Line 16   Column 84   Coefficient 0.00001144
         when "111101010100" => A <= "000000000000000100"; -- Line 16   Column 85   Coefficient 0.00001526
         when "111101010101" => A <= "000000000000000110"; -- Line 16   Column 86   Coefficient 0.00002289
         when "111101010110" => A <= "000000000000000011"; -- Line 16   Column 87   Coefficient 0.00001144
         when "111101010111" => A <= "111111111111111111"; -- Line 16   Column 88   Coefficient -0.00000381
         when "111101011000" => A <= "000000000000000000"; -- Line 16   Column 89   Coefficient 0.00000000
         when "111101011001" => A <= "000000000000000000"; -- Line 16   Column 90   Coefficient 0.00000000
         when "111101011010" => A <= "000000000000000000"; -- Line 16   Column 91   Coefficient 0.00000000
         when "111101011011" => A <= "000000000000000000"; -- Line 16   Column 92   Coefficient 0.00000000
         when "111101011100" => A <= "000000000000000000"; -- Line 16   Column 93   Coefficient 0.00000000
         when "111101011101" => A <= "000000000000000000"; -- Line 16   Column 94   Coefficient 0.00000000
         when "111101011110" => A <= "000000000000000000"; -- Line 16   Column 95   Coefficient 0.00000000
         when "111101011111" => A <= "000000000000000000"; -- Line 16   Column 96   Coefficient 0.00000000
         when "111101100000" => A <= "000000000000000000"; -- Line 16   Column 97   Coefficient 0.00000000
         when "111101100001" => A <= "000000000000000000"; -- Line 16   Column 98   Coefficient 0.00000000
         when "111101100010" => A <= "000000000000000000"; -- Line 16   Column 99   Coefficient 0.00000000
         when "111101100011" => A <= "000000000000000000"; -- Line 16   Column 100   Coefficient 0.00000000
         when "111101100100" => A <= "000000000000000000"; -- Line 16   Column 101   Coefficient 0.00000000
         when "111101100101" => A <= "000000000000000000"; -- Line 16   Column 102   Coefficient 0.00000000
         when "111101100110" => A <= "000000000000000000"; -- Line 16   Column 103   Coefficient 0.00000000
         when "111101100111" => A <= "000000000000000000"; -- Line 16   Column 104   Coefficient 0.00000000
         when "111101101000" => A <= "000000000000000000"; -- Line 16   Column 105   Coefficient 0.00000000
         when "111101101001" => A <= "000000000000000000"; -- Line 16   Column 106   Coefficient 0.00000000
         when "111101101010" => A <= "000000000000000000"; -- Line 16   Column 107   Coefficient 0.00000000
         when "111101101011" => A <= "000000000000000000"; -- Line 16   Column 108   Coefficient 0.00000000
         when "111101101100" => A <= "000000000000000000"; -- Line 16   Column 109   Coefficient 0.00000000
         when "111101101101" => A <= "000000000000000000"; -- Line 16   Column 110   Coefficient 0.00000000
         when "111101101110" => A <= "000000000000000000"; -- Line 16   Column 111   Coefficient 0.00000000
         when "111101101111" => A <= "000000000000000000"; -- Line 16   Column 112   Coefficient 0.00000000
         when "111101110000" => A <= "000000000000000000"; -- Line 16   Column 113   Coefficient 0.00000000
         when "111101110001" => A <= "000000000000000000"; -- Line 16   Column 114   Coefficient 0.00000000
         when "111101110010" => A <= "000000000000000000"; -- Line 16   Column 115   Coefficient 0.00000000
         when "111101110011" => A <= "000000000000000000"; -- Line 16   Column 116   Coefficient 0.00000000
         when "111101110100" => A <= "000000000000000000"; -- Line 16   Column 117   Coefficient 0.00000000
         when "111101110101" => A <= "000000000000000000"; -- Line 16   Column 118   Coefficient 0.00000000
         when "111101110110" => A <= "000000000000000000"; -- Line 16   Column 119   Coefficient 0.00000000
         when "111101110111" => A <= "000000000000000000"; -- Line 16   Column 120   Coefficient 0.00000000
         when "111101111000" => A <= "000000000000000000"; -- Line 16   Column 121   Coefficient 0.00000000
         when "111101111001" => A <= "000000000000000000"; -- Line 16   Column 122   Coefficient 0.00000000
         when "111101111010" => A <= "000000000000000000"; -- Line 16   Column 123   Coefficient 0.00000000
         when "111101111011" => A <= "000000000000000000"; -- Line 16   Column 124   Coefficient 0.00000000
         when "111101111100" => A <= "000000000000000000"; -- Line 16   Column 125   Coefficient 0.00000000
         when "111101111101" => A <= "000000000000000000"; -- Line 16   Column 126   Coefficient 0.00000000
         when "111101111110" => A <= "000000000000000000"; -- Line 16   Column 127   Coefficient 0.00000000
         when "111101111111" => A <= "000000000000000000"; -- Line 16   Column 128   Coefficient 0.00000000
         when "111110000000" => A <= "000000000000000000"; -- Line 16   Column 129   Coefficient 0.00000000
         when "111110000001" => A <= "000000000000000000"; -- Line 16   Column 130   Coefficient 0.00000000
         when "111110000010" => A <= "000000000000000000"; -- Line 16   Column 131   Coefficient 0.00000000
         when "111110000011" => A <= "000000000000000000"; -- Line 16   Column 132   Coefficient 0.00000000
         when "111110000100" => A <= "000000000000000000"; -- Line 16   Column 133   Coefficient 0.00000000
         when "111110000101" => A <= "000000000000000000"; -- Line 16   Column 134   Coefficient 0.00000000
         when "111110000110" => A <= "000000000000000000"; -- Line 16   Column 135   Coefficient 0.00000000
         when "111110000111" => A <= "000000000000000000"; -- Line 16   Column 136   Coefficient 0.00000000
         when "111110001000" => A <= "000000000000000000"; -- Line 16   Column 137   Coefficient 0.00000000
         when "111110001001" => A <= "000000000000000000"; -- Line 16   Column 138   Coefficient 0.00000000
         when "111110001010" => A <= "000000000000000000"; -- Line 16   Column 139   Coefficient 0.00000000
         when "111110001011" => A <= "000000000000000000"; -- Line 16   Column 140   Coefficient 0.00000000
         when "111110001100" => A <= "000000000000000000"; -- Line 16   Column 141   Coefficient 0.00000000
         when "111110001101" => A <= "000000000000000000"; -- Line 16   Column 142   Coefficient 0.00000000
         when "111110001110" => A <= "000000000000000000"; -- Line 16   Column 143   Coefficient 0.00000000
         when "111110001111" => A <= "000000000000000000"; -- Line 16   Column 144   Coefficient 0.00000000
         when "111110010000" => A <= "000000000000000000"; -- Line 16   Column 145   Coefficient 0.00000000
         when "111110010001" => A <= "000000000000000000"; -- Line 16   Column 146   Coefficient 0.00000000
         when "111110010010" => A <= "000000000000000000"; -- Line 16   Column 147   Coefficient 0.00000000
         when "111110010011" => A <= "000000000000000000"; -- Line 16   Column 148   Coefficient 0.00000000
         when "111110010100" => A <= "000000000000000000"; -- Line 16   Column 149   Coefficient 0.00000000
         when "111110010101" => A <= "000000000000000000"; -- Line 16   Column 150   Coefficient 0.00000000
         when "111110010110" => A <= "000000000000000000"; -- Line 16   Column 151   Coefficient 0.00000000
         when "111110010111" => A <= "000000000000000000"; -- Line 16   Column 152   Coefficient 0.00000000
         when "111110011000" => A <= "000000000000000000"; -- Line 16   Column 153   Coefficient 0.00000000
         when "111110011001" => A <= "000000000000000000"; -- Line 16   Column 154   Coefficient 0.00000000
         when "111110011010" => A <= "000000000000000000"; -- Line 16   Column 155   Coefficient 0.00000000
         when "111110011011" => A <= "000000000000000000"; -- Line 16   Column 156   Coefficient 0.00000000
         when "111110011100" => A <= "000000000000000000"; -- Line 16   Column 157   Coefficient 0.00000000
         when "111110011101" => A <= "000000000000000000"; -- Line 16   Column 158   Coefficient 0.00000000
         when "111110011110" => A <= "000000000000000000"; -- Line 16   Column 159   Coefficient 0.00000000
         when "111110011111" => A <= "000000000000000000"; -- Line 16   Column 160   Coefficient 0.00000000
         when "111110100000" => A <= "000000000000000000"; -- Line 16   Column 161   Coefficient 0.00000000
         when "111110100001" => A <= "000000000000000000"; -- Line 16   Column 162   Coefficient 0.00000000
         when "111110100010" => A <= "000000000000000000"; -- Line 16   Column 163   Coefficient 0.00000000
         when "111110100011" => A <= "000000000000000000"; -- Line 16   Column 164   Coefficient 0.00000000
         when "111110100100" => A <= "000000000000000000"; -- Line 16   Column 165   Coefficient 0.00000000
         when "111110100101" => A <= "000000000000000000"; -- Line 16   Column 166   Coefficient 0.00000000
         when "111110100110" => A <= "000000000000000000"; -- Line 16   Column 167   Coefficient 0.00000000
         when "111110100111" => A <= "000000000000000000"; -- Line 16   Column 168   Coefficient 0.00000000
         when "111110101000" => A <= "000000000000000000"; -- Line 16   Column 169   Coefficient 0.00000000
         when "111110101001" => A <= "000000000000000000"; -- Line 16   Column 170   Coefficient 0.00000000
         when "111110101010" => A <= "000000000000000000"; -- Line 16   Column 171   Coefficient 0.00000000
         when "111110101011" => A <= "000000000000000000"; -- Line 16   Column 172   Coefficient 0.00000000
         when "111110101100" => A <= "000000000000000000"; -- Line 16   Column 173   Coefficient 0.00000000
         when "111110101101" => A <= "000000000000000000"; -- Line 16   Column 174   Coefficient 0.00000000
         when "111110101110" => A <= "000000000000000000"; -- Line 16   Column 175   Coefficient 0.00000000
         when "111110101111" => A <= "000000000000000000"; -- Line 16   Column 176   Coefficient 0.00000000
         when "111110110000" => A <= "000000000000000000"; -- Line 16   Column 177   Coefficient 0.00000000
         when "111110110001" => A <= "000000000000000000"; -- Line 16   Column 178   Coefficient 0.00000000
         when "111110110010" => A <= "000000000000000000"; -- Line 16   Column 179   Coefficient 0.00000000
         when "111110110011" => A <= "000000000000000000"; -- Line 16   Column 180   Coefficient 0.00000000
         when "111110110100" => A <= "000000000000000000"; -- Line 16   Column 181   Coefficient 0.00000000
         when "111110110101" => A <= "000000000000000000"; -- Line 16   Column 182   Coefficient 0.00000000
         when "111110110110" => A <= "000000000000000000"; -- Line 16   Column 183   Coefficient 0.00000000
         when "111110110111" => A <= "000000000000000000"; -- Line 16   Column 184   Coefficient 0.00000000
         when "111110111000" => A <= "000000000000000000"; -- Line 16   Column 185   Coefficient 0.00000000
         when "111110111001" => A <= "000000000000000000"; -- Line 16   Column 186   Coefficient 0.00000000
         when "111110111010" => A <= "000000000000000000"; -- Line 16   Column 187   Coefficient 0.00000000
         when "111110111011" => A <= "000000000000000000"; -- Line 16   Column 188   Coefficient 0.00000000
         when "111110111100" => A <= "000000000000000000"; -- Line 16   Column 189   Coefficient 0.00000000
         when "111110111101" => A <= "000000000000000000"; -- Line 16   Column 190   Coefficient 0.00000000
         when "111110111110" => A <= "000000000000000000"; -- Line 16   Column 191   Coefficient 0.00000000
         when "111110111111" => A <= "000000000000000000"; -- Line 16   Column 192   Coefficient 0.00000000
         when "111111000000" => A <= "000000000000000000"; -- Line 16   Column 193   Coefficient 0.00000000
         when "111111000001" => A <= "000000000000000000"; -- Line 16   Column 194   Coefficient 0.00000000
         when "111111000010" => A <= "000000000000000000"; -- Line 16   Column 195   Coefficient 0.00000000
         when "111111000011" => A <= "000000000000000000"; -- Line 16   Column 196   Coefficient 0.00000000
         when "111111000100" => A <= "000000000000000000"; -- Line 16   Column 197   Coefficient 0.00000000
         when "111111000101" => A <= "000000000000000000"; -- Line 16   Column 198   Coefficient 0.00000000
         when "111111000110" => A <= "000000000000000000"; -- Line 16   Column 199   Coefficient 0.00000000
         when "111111000111" => A <= "000000000000000000"; -- Line 16   Column 200   Coefficient 0.00000000
         when "111111001000" => A <= "000000000000000000"; -- Line 16   Column 201   Coefficient 0.00000000
         when "111111001001" => A <= "000000000000000000"; -- Line 16   Column 202   Coefficient 0.00000000
         when "111111001010" => A <= "000000000000000000"; -- Line 16   Column 203   Coefficient 0.00000000
         when "111111001011" => A <= "000000000000000000"; -- Line 16   Column 204   Coefficient 0.00000000
         when "111111001100" => A <= "000000000000000000"; -- Line 16   Column 205   Coefficient 0.00000000
         when "111111001101" => A <= "000000000000000000"; -- Line 16   Column 206   Coefficient 0.00000000
         when "111111001110" => A <= "000000000000000000"; -- Line 16   Column 207   Coefficient 0.00000000
         when "111111001111" => A <= "000000000000000000"; -- Line 16   Column 208   Coefficient 0.00000000
         when "111111010000" => A <= "000000000000000000"; -- Line 16   Column 209   Coefficient 0.00000000
         when "111111010001" => A <= "000000000000000000"; -- Line 16   Column 210   Coefficient 0.00000000
         when "111111010010" => A <= "000000000000000000"; -- Line 16   Column 211   Coefficient 0.00000000
         when "111111010011" => A <= "000000000000000000"; -- Line 16   Column 212   Coefficient 0.00000000
         when "111111010100" => A <= "000000000000000000"; -- Line 16   Column 213   Coefficient 0.00000000
         when "111111010101" => A <= "000000000000000000"; -- Line 16   Column 214   Coefficient 0.00000000
         when "111111010110" => A <= "000000000000000000"; -- Line 16   Column 215   Coefficient 0.00000000
         when "111111010111" => A <= "000000000000000000"; -- Line 16   Column 216   Coefficient 0.00000000
         when "111111011000" => A <= "000000000000000000"; -- Line 16   Column 217   Coefficient 0.00000000
         when "111111011001" => A <= "000000000000000000"; -- Line 16   Column 218   Coefficient 0.00000000
         when "111111011010" => A <= "000000000000000000"; -- Line 16   Column 219   Coefficient 0.00000000
         when "111111011011" => A <= "000000000000000000"; -- Line 16   Column 220   Coefficient 0.00000000
         when "111111011100" => A <= "000000000000000000"; -- Line 16   Column 221   Coefficient 0.00000000
         when "111111011101" => A <= "000000000000000000"; -- Line 16   Column 222   Coefficient 0.00000000
         when "111111011110" => A <= "000000000000000000"; -- Line 16   Column 223   Coefficient 0.00000000
         when "111111011111" => A <= "000000000000000000"; -- Line 16   Column 224   Coefficient 0.00000000
         when "111111100000" => A <= "000000000000000000"; -- Line 16   Column 225   Coefficient 0.00000000
         when "111111100001" => A <= "000000000000000000"; -- Line 16   Column 226   Coefficient 0.00000000
         when "111111100010" => A <= "000000000000000000"; -- Line 16   Column 227   Coefficient 0.00000000
         when "111111100011" => A <= "000000000000000000"; -- Line 16   Column 228   Coefficient 0.00000000
         when "111111100100" => A <= "000000000000000000"; -- Line 16   Column 229   Coefficient 0.00000000
         when "111111100101" => A <= "000000000000000000"; -- Line 16   Column 230   Coefficient 0.00000000
         when "111111100110" => A <= "000000000000000000"; -- Line 16   Column 231   Coefficient 0.00000000
         when "111111100111" => A <= "000000000000000000"; -- Line 16   Column 232   Coefficient 0.00000000
         when "111111101000" => A <= "000000000000000000"; -- Line 16   Column 233   Coefficient 0.00000000
         when "111111101001" => A <= "000000000000000000"; -- Line 16   Column 234   Coefficient 0.00000000
         when "111111101010" => A <= "000000000000000000"; -- Line 16   Column 235   Coefficient 0.00000000
         when "111111101011" => A <= "000000000000000000"; -- Line 16   Column 236   Coefficient 0.00000000
         when "111111101100" => A <= "000000000000000000"; -- Line 16   Column 237   Coefficient 0.00000000
         when "111111101101" => A <= "000000000000000000"; -- Line 16   Column 238   Coefficient 0.00000000
         when "111111101110" => A <= "000000000000000000"; -- Line 16   Column 239   Coefficient 0.00000000
         when "111111101111" => A <= "000000000000000000"; -- Line 16   Column 240   Coefficient 0.00000000
         when "111111110000" => A <= "000000000000001001"; -- Line 16   Column 241   Coefficient 0.00003433
         when "111111110001" => A <= "000000000000000011"; -- Line 16   Column 242   Coefficient 0.00001144
         when "111111110010" => A <= "111111111111001011"; -- Line 16   Column 243   Coefficient -0.00020218
         when "111111110011" => A <= "111111111110100110"; -- Line 16   Column 244   Coefficient -0.00034332
         when "111111110100" => A <= "111111111110010010"; -- Line 16   Column 245   Coefficient -0.00041962
         when "111111110101" => A <= "111111111111010011"; -- Line 16   Column 246   Coefficient -0.00017166
         when "111111110110" => A <= "000000000011111000"; -- Line 16   Column 247   Coefficient 0.00094604
         when "111111110111" => A <= "000000001000010011"; -- Line 16   Column 248   Coefficient 0.00202560
         when "111111111000" => A <= "000000001010110110"; -- Line 16   Column 249   Coefficient 0.00264740
         when "111111111001" => A <= "000000001101001100"; -- Line 16   Column 250   Coefficient 0.00321960
         when "111111111010" => A <= "000000001111111100"; -- Line 16   Column 251   Coefficient 0.00389099
         when "111111111011" => A <= "000000010000011000"; -- Line 16   Column 252   Coefficient 0.00399780
         when "111111111100" => A <= "000000001111000010"; -- Line 16   Column 253   Coefficient 0.00366974
         when "111111111101" => A <= "000000000111011010"; -- Line 16   Column 254   Coefficient 0.00180817
         when "111111111110" => A <= "111111110001010101"; -- Line 16   Column 255   Coefficient -0.00358200
         when "111111111111" => A <= "111111011001111001"; -- Line 16   Column 256   Coefficient -0.00930405
         when others => null;
      end case;
   end process;
end LUTable;
